// Verilog netlist created by TD v4.6.18154
// Thu Nov 12 15:31:47 2020

`timescale 1ns / 1ps
module rom_wb1  // al_ip/ann/rom_wb1.v(14)
  (
  addra,
  clka,
  rsta,
  doa
  );

  input [9:0] addra;  // al_ip/ann/rom_wb1.v(18)
  input clka;  // al_ip/ann/rom_wb1.v(19)
  input rsta;  // al_ip/ann/rom_wb1.v(20)
  output [449:0] doa;  // al_ip/ann/rom_wb1.v(16)


  EG_PHY_CONFIG #(
    .DONE_PERSISTN("ENABLE"),
    .INIT_PERSISTN("ENABLE"),
    .JTAG_PERSISTN("DISABLE"),
    .PROGRAMN_PERSISTN("DISABLE"))
    config_inst ();
  // address_offset=0;data_offset=0;depth=785;width=9;num_section=1;width_per_section=9;section_size=450;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hA467FC8262051C1083878A11D8C33031F8D242EC1E1781A17E3FE7EED64F2710),
    .INITP_01(256'hE0A501FE62A83FEC0FF7FEC2677940307E001387C00320100071FC85181F8F14),
    .INITP_02(256'h407BCBBCF97E818687C6053414484189806A9DBB0E36087680E19F815F074817),
    .INITP_03(256'h000000000000000000000000000000000000000000000000000000000000E8BB),
    .INIT_00(256'h0C06000708070B01030200050303040100090400050404050009050106070016),
    .INIT_01(256'h02020706020B0900050001140A15100714201429650A32330F0F11000B070108),
    .INIT_02(256'h30581B020C6A040E21010001000117151A3C2A1652430E142C0C392319010023),
    .INIT_03(256'h13633A312A1A1A10160825072F0401061C13364F384D13041D210E107920090D),
    .INIT_04(256'h07040A2D05081F130609151729360452180E020159264A5E24340307243D1007),
    .INIT_05(256'h1E011C122119110A0801000F070C2516102C2A08100C010E333441030D29060E),
    .INIT_06(256'h5E3B1C01150B151822050A1206050014110300024B240E15075200073A271418),
    .INIT_07(256'h1927023F0843230704010E090901180C1702191701051B2A0D06312F0D4B650B),
    .INIT_08(256'h12083F3311250B137F1114020E03454E1E010E0D100C3010060B1C09000F3B1B),
    .INIT_09(256'h252300171B12572F013B0122330C1E1B1E021C29120F0001140E0A1C2E011306),
    .INIT_0A(256'h26182624121024510A203C53450D011E360D151D0303060912071409012C532E),
    .INIT_0B(256'h04093B3221431A1E19151C1907210050600700060615130313080B0F03140A1C),
    .INIT_0C(256'h0C08200006103C40081B551C0709291D0D02017B3606190A6A2617052523000E),
    .INIT_0D(256'h2D1C021306221203162807072B01403D4B1D17290E3F3F580A180E0444212A1C),
    .INIT_0E(256'h0004031332092C1C20040E0705001E153C1434665B284149162261470411040D),
    .INIT_0F(256'h21160C191902471F130D0906170222030D0C211D331909081C26246B2C2D5124),
    .INIT_10(256'h110117151A3F4D0C695E073A330A222C0F0425020409052A323B16170819325A),
    .INIT_11(256'h060A020F230E2501041B5A253C00000901280D111D221D05130016112C3A200A),
    .INIT_12(256'h0D220C160E030912191E0B0B1E01213C060B02070A26180C0019141504060425),
    .INIT_13(256'h030B0B0015200A0D110F070F0B0C021306183C083C0205016C2920051A1F1B02),
    .INIT_14(256'h0A52070601112D1F03071B1A14150B020F080401092F5E22140103004751031E),
    .INIT_15(256'h2E00050200385D5F472B02461935100E04052F220B0F0A1E18073D3A0C020008),
    .INIT_16(256'h383D4E0301000405021D0B57390E19140201072C20071D2439140B002837263B),
    .INIT_17(256'h06082823151F0E05000804050A0717261810131B06001A3327272F2346131607),
    .INIT_18(256'h000000000000000000000000000000030703010914024B13353422364F02020A),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_785x450_sub_000000_000 (
    .addra({addra,3'b111}),
    .clka(clka),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa(doa[8:0]));
  // address_offset=0;data_offset=9;depth=785;width=9;num_section=1;width_per_section=9;section_size=450;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h49C1FBCD1FAFDBF4FD91783C9864505006E0DC67C0D0FFFFF46F9FF0B57CFDF9),
    .INITP_01(256'h02EA1FEC10371FE341C1FE1CF009F93E003FF783037FFE580FFC81F067181F0E),
    .INITP_02(256'hFE4706E6F840BD3F2E3C08429F000F3F4827C3EC2EE0FE81FC0F6C1F40FEE9FC),
    .INITP_03(256'h000000000000000000000000000000000000000000000000000000000001574F),
    .INIT_00(256'h05000D03010D0901040101030902000006020305020705020105010703000406),
    .INIT_01(256'h0B0A080B0004010A0701020305040D05070A0D09030B1B0A0B18070F03000002),
    .INIT_02(256'h3E47420D3A3E1C070B07040404050D060C242A3934438D776E8B4B3C0732060C),
    .INIT_03(256'h1D041D2734010D09021E1F4D0D080007084415222A1C34070B1106022203354B),
    .INIT_04(256'h1C1A082004131B180808283421330A26310307073D1F581A051F01081F1E3944),
    .INIT_05(256'h0E19040F1E030401011004040C0A0F1A11121F41150E020F1C15071A1D2A0C0E),
    .INIT_06(256'h4A43183A0A160F04060E04100F140C190604112A0A320E1E2A4301014C1B1D0A),
    .INIT_07(256'h372103130565124105181B18201C011905171E150421061D3B1A032F015E0105),
    .INIT_08(256'h0E2F65002B18060D0647070B0B08181A10091B19191E0A0C04151A061338480D),
    .INIT_09(256'h07080A1405486A3935160B30441C161506091316110A0510060E06301110291A),
    .INIT_0A(256'h0D1C40303B0616280339804220050B342A1F2E1A42160C14150F1F0A05044105),
    .INIT_0B(256'h170A06172B37452D072013300B3635242712031B340B3E3C2D1D050811000210),
    .INIT_0C(256'h4F431A180F210F21394C340B1D030F24302E641C3F03090C061E221E35150E00),
    .INIT_0D(256'h3A071A2C1D00041C21050F0C22393706293F1D43285214022F1003160D0B071A),
    .INIT_0E(256'h2D070002214A1A0E261A2516070A0404000A15226252343B256A0A3242150A0A),
    .INIT_0F(256'h47445A44180A590B423D122D06281B0003070F1B170E332B640B020E04023C12),
    .INIT_10(256'h010A0C2530561C7D04600A2C645308271C24043A010C1601372D55122F052642),
    .INIT_11(256'h0C121101021A00140F2A315C1F06012414350D1B1E090E26330B271C353C440E),
    .INIT_12(256'h0F17060A0E1827052E2A1A04181D16112B111008075D09260910261525131E09),
    .INIT_13(256'h1B1005200209010205071117063232200715241302020907133D5003160B1118),
    .INIT_14(256'h25262F291F14222D0006060C1D19072D25142636070926092806080204184113),
    .INIT_15(256'h19000C02160B1D01282D04320D152E1B1D0E320D02272D40291F0A1C01010208),
    .INIT_16(256'h30822116020213040C082E403B36290B1E000A0A020917241B1408241E030614),
    .INIT_17(256'h492B2D20160A07020002010F04070245293C2A130B06090413632A141A092017),
    .INIT_18(256'h000000000000000000000000000000080B01000708234C082349001C23123C3A),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_785x450_sub_000000_009 (
    .addra({addra,3'b111}),
    .clka(clka),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa(doa[17:9]));
  // address_offset=0;data_offset=18;depth=785;width=9;num_section=1;width_per_section=9;section_size=450;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFE007004E00703CCCFF81E8CF7068800609DC31E01B223E03E597013E24184D2),
    .INITP_01(256'hE71106505A801D2F66B8C259634839A7CF863D3DD821DBFC00196FF09388CF02),
    .INITP_02(256'h38D3FBFFD6C32ABC8EC5BFFBA013BC70A813DA2B001C5FE006F1D947BED59C19),
    .INITP_03(256'h000000000000000000000000000000000000000000000000000000000000F9F2),
    .INIT_00(256'h090404020109070209040400040105050305090206040005060309010402021F),
    .INIT_01(256'h0F060D1F01080102000400060A08100B20011B0A2C13212D2B1B0B0602050202),
    .INIT_02(256'h242F081300162018240E04090302041F4409021D321E222108122C070735271B),
    .INIT_03(256'h013B2424393E201225041129300102011C05368A15022F05010802132E6B2B2D),
    .INIT_04(256'h010F0E0F124A44111F26171E0C175F0D1B05003313203F442422191C0D122D1A),
    .INIT_05(256'h0B1426251B030B0A122C322E24211F0B22461C141A08093225032A0C12050F1E),
    .INIT_06(256'h0A792C203C230C1603141B20072F3A28062222110E431F04081100252D190B1A),
    .INIT_07(256'h160A011D0A2C0A030A230B0D100B190D0C1E3D1B10313F3339302C0913055B2B),
    .INIT_08(256'h0F11162F0E0503301F381409171D0A12060B08080532491C0E2D2B291E050E04),
    .INIT_09(256'h1E2F211F3221051A290704245E283A150D120C0017171314252C211D182B110E),
    .INIT_0A(256'h4C05130D091228370C00193F32020728342602201E02232D38291616283B1001),
    .INIT_0B(256'h171E020F110F0414191513280D090A230912042B1306361B020A2D322110100A),
    .INIT_0C(256'h1E0F2210070E08030015140A1D090A22232F26210F000A02720508111D022725),
    .INIT_0D(256'h1B10153A14150B0705170410010411210E160A2D180304132A0111083D010707),
    .INIT_0E(256'h300204350E0D13120100091104122A22010214041E0C1202000E0A4211050433),
    .INIT_0F(256'h180C073B2D0A2638422E180E1505150C140431210B05040D1105030E060A061E),
    .INIT_10(256'h0D04051316191E4126060C3A2B0C1A1C12080D150E190B0E15150C2B0803001D),
    .INIT_11(256'h14171C1018050800172A4F070E08002A09162A160900000D000B00171F170812),
    .INIT_12(256'h071C0A1A25371F030903011728520819040701041026170802090F0031091324),
    .INIT_13(256'h0712081407112C24181318150C070A1B46173C203B0507001B0027220403071F),
    .INIT_14(256'h14121E0F152514261F090812090112390209394E0C101D1F040A01091400020B),
    .INIT_15(256'h2B0A0204101328020B0923021A180F1706090D06221B72364D3F030521000507),
    .INIT_16(256'h58470005000405000E143A5B2D13141D26020F130A1D0B0C32100A263450180D),
    .INIT_17(256'h27001C15140A06070209040700041A0D55257145120021444628150B35033D58),
    .INIT_18(256'h000000000000000000000000000000000106020820284C48400E42270045231E),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_785x450_sub_000000_018 (
    .addra({addra,3'b111}),
    .clka(clka),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa(doa[26:18]));
  // address_offset=0;data_offset=27;depth=785;width=9;num_section=1;width_per_section=9;section_size=450;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h2F740034FFC221077800037A380421FFC3E71FFFC06D3DCFCA4147022CA98DE5),
    .INITP_01(256'h8840F8789C3F819B83E401B8BE00E3ABAACEF320FDC5041F941C01F94F882100),
    .INITP_02(256'h00600000228809033E540001A400FB5B405F17F01E612407EDD0407DD9360FC7),
    .INITP_03(256'h000000000000000000000000000000000000000000000000000000000000A300),
    .INIT_00(256'h040302090301040403020D0505000B01050B0805030202030203080001010730),
    .INIT_01(256'h110210080100080004010504050C0201010811090D02070D0903070304050605),
    .INIT_02(256'h07404C39385A080E070507010B0902061411314850090B16574F2035062C3104),
    .INIT_03(256'h303D16292519192F1F3D12581106070100021113211B3B525016274845353101),
    .INIT_04(256'h2A08081C1400094E24482B18151B19090A090501060D1E184B01284E1C373424),
    .INIT_05(256'h080724152103043914211B323616072C061312142E0C03042A1220650C000C15),
    .INIT_06(256'h2A6548421719151201230F3F283D05150E00040F3A130A2E3B0F00203C0C585D),
    .INIT_07(256'h06000416244F143108190F050A061604133731150D102A0A3710100F18040D27),
    .INIT_08(256'h180A28481006013A1E141C0B0E092800162901040F0B1214062D111610071B28),
    .INIT_09(256'h17070714001008490F11004A031A033424185204261D150A02092124141C0D09),
    .INIT_0A(256'h1A1F360C3102040C030E281C0001023B3853380B0B081E342228161026100610),
    .INIT_0B(256'h1A01040C03072303051A0E0510140908020C1023052031021C182707191E0A00),
    .INIT_0C(256'h1106154319022403031A02241C0D08000B2E1D0A130D08141A0E06090C250F2C),
    .INIT_0D(256'h580D6E3528100B1706041D0600040A2E2D0D1B09040D031F32120217661A3424),
    .INIT_0E(256'h3D0500213023382E3507121921251B111D020417220001031615261637170602),
    .INIT_0F(256'h061D131C370F440D0129083C17030B0033232C1E05010103040E190B221D2C2E),
    .INIT_10(256'h370F0F190E1B0C130C160613613A161830244437101835161F16060C0C01070B),
    .INIT_11(256'h0E330101050A0B153A18051B00100906496D10074F2936500806100413302D0C),
    .INIT_12(256'h1005090711330F040D382E0E1E1D2C1B3B0F0804101D0C072D2A233D2016091B),
    .INIT_13(256'h15070E0F1E36211D0B19051F162E441A070E1A34010105060A0514121C0A171F),
    .INIT_14(256'h4A072F00121F060420132248272D1117030F1D091C10141039050A073B003A16),
    .INIT_15(256'h3504010734650432190300170C18051417514925251326343318123B1B070401),
    .INIT_16(256'h603705070003030002004D010B0E1C4C111410081A102602442F472F08210C15),
    .INIT_17(256'h1507201C0B00030301030A09000118565C278F667B402E2F7A77535D301D5475),
    .INIT_18(256'h0000000000000000000000000000000401060B1D573A3411616D4C23573C503D),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_785x450_sub_000000_027 (
    .addra({addra,3'b111}),
    .clka(clka),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa(doa[35:27]));
  // address_offset=0;data_offset=36;depth=785;width=9;num_section=1;width_per_section=9;section_size=450;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h5990617600089E441001D577B03F9732FF8ED13FFF97FFFFF47FF8FE0301738C),
    .INITP_01(256'h743F0E076BD3C5DF7F3E5CFB46849BB06809BF86E0077A060369E77016950407),
    .INITP_02(256'h07CC100A0BB1960E5E5F20F183F147E9FD723C99EFFBE941DFB9301DCDF7E86C),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000001C44),
    .INIT_00(256'h07020005040A02080005020700040504000415030300050301020A010604022A),
    .INIT_01(256'h1204333900050902010404342923441F232F2D330E09140D1A1E211615080702),
    .INIT_02(256'h58540E1D2115444202000003000A2D48395B38410A1C7B786E799E824F312A0C),
    .INIT_03(256'h3339595A44767D1411040103020601000502073508141D0E1B0A2428798F442B),
    .INIT_04(256'h200239210C1E1A18251615613D012C0816050218001511044D141B350A261408),
    .INIT_05(256'h32381612062D05070D00220F08371E36582520012D0F05121625404107091637),
    .INIT_06(256'h7A12293729060D2820431815010E07000515165E283E090234260C01741D0321),
    .INIT_07(256'h08030022357E371A0F01042926191C2D2F111217070A4832113E050E231F3204),
    .INIT_08(256'h181B10021317091D532F33390108122B010A0A062D09090B0E052D120C062316),
    .INIT_09(256'h2424372C0F092C1A477302133E1A1E4205101B0E060812021F202108031D232B),
    .INIT_0A(256'h13161F1324164111020E2F0253090418111F0E39090618011C0E100104230709),
    .INIT_0B(256'h052C0806013019042A082D260C1A260C2101180C1C1330100E05001715120B04),
    .INIT_0C(256'h3907181A27080E001025160E0A060D2614020E262D0011305F2E3D0E1B010806),
    .INIT_0D(256'h1E1243190216020616131D0E1A0101120515111912194D0201080C06200E440B),
    .INIT_0E(256'h0413020706064810223714090328160A2008161A021C12391D1B151B0F200A02),
    .INIT_0F(256'h031D0F08160B141030303A4A1D40081B0A26170D0A0809092E2A0F0010183615),
    .INIT_10(256'h363C0B130D0C0303031801443437703418332C00101B240F051A19020F030E0B),
    .INIT_11(256'h02211C0D3E460430060014270E50052C0A294924000A0220230B020C101C1F25),
    .INIT_12(256'h1702030E15390C24472B1E21253D01184A1B03032E6D1D1314051F230308170A),
    .INIT_13(256'h1F1206112C130910062C222A0A12030D1D0545194B0300006F2E2511240E060E),
    .INIT_14(256'h085827311206120E0E011A1A0E00020307090A081B266A1443050706244F2A04),
    .INIT_15(256'h1C02070D08231F372F0A13071B352304091C011F1B0B1925031E132001000205),
    .INIT_16(256'h2E446213010006060B09511810110E0D180C0F0F00233A141615302F2606110A),
    .INIT_17(256'h100B1B211C17040104060001040C2A49452E102E030C080239071D0204180321),
    .INIT_18(256'h0000000000000000000000000000000D07010518130803531946001D0408221F),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_785x450_sub_000000_036 (
    .addra({addra,3'b111}),
    .clka(clka),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa(doa[44:36]));
  // address_offset=0;data_offset=45;depth=785;width=9;num_section=1;width_per_section=9;section_size=450;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h08476043983A061F004001BF10DB30B0FFC083DFFB83FBFFFC3FF3FBE081C50A),
    .INITP_01(256'h3833A3B4F4003EC83C02F4A3CE06023903182382E582303C04410F2E0220E482),
    .INITP_02(256'h780B0010EC3F8668ECFFEC11DFFEE5DCFDD017DF99D938FBBFE7FB93B127B837),
    .INITP_03(256'h000000000000000000000000000000000000000000000000000000000001C100),
    .INIT_00(256'h0B02060000050508050002040306060302010607060503030300060103070420),
    .INIT_01(256'h0C092F43090402040700081D20203A2A272819301B0513070C20151203010A04),
    .INIT_02(256'h3E9A6A65380A314C0A04010904000F22435E34450D18134E47249F7F6C1A110B),
    .INIT_03(256'h0F223F4130B04617220F2C0F12030E041E0F2C3A0F1F35573B20140138A1630C),
    .INIT_04(256'h35371B0E00122B200A01411C29070739040404210F272907040E021122250006),
    .INIT_05(256'h1836120E2335170C0F1A2006244606090530334C170803250627023E1C0A1218),
    .INIT_06(256'h44304403050C2C2027220F081205040E0000001C1B2C0E906059022E010F0705),
    .INIT_07(256'h1B4C00030A2911160B1424181D14270F15101E0A0E062612112B1C4459616023),
    .INIT_08(256'h1E1F152B3A0401495321060B192E551F0F124D01200214110C15000A0B20023E),
    .INIT_09(256'h290C121A0C0602323D4F01655E0300250F3D490F03052C2207140A0606061318),
    .INIT_0A(256'h023316062D06020E02341A175C1202542B0533351C1B200D00062C22030C1426),
    .INIT_0B(256'h0E0113020C0403081D010310062D261D64111C56430441572C211D24250F0B0D),
    .INIT_0C(256'h27060E221006070B0A3128180619051A120026102E11101A3A33265C26343803),
    .INIT_0D(256'h093342220B200C1303040D2C1C10060B071A23110C2F132C47000B0F160C4D24),
    .INIT_0E(256'h280C01103346040F002012020419050A1E151C45050C2102032007115A0D0610),
    .INIT_0F(256'h040517030407470B2F133B05160D071B0918041C192623351718050903210E0F),
    .INIT_10(256'h13100628030C011E3B4E10004C0955691F1D23031C1814020414210E00281B11),
    .INIT_11(256'h05261D06140204270C0B492326290A391B1B2F2A2E002E04250D0815081E1323),
    .INIT_12(256'h1C230820261812040E0204290E2E21211A1D18030E4F3E2321181C172D011211),
    .INIT_13(256'h0637412C09040B24271605090A0B2C191519151B3B0A19076E281E11221D310C),
    .INIT_14(256'h530A0F1104432527160111183B241808030C081B211A005B3605060466291C06),
    .INIT_15(256'h1C160100263B0B0003330D1F1E0104170C2E360A082108192026153C22000D0A),
    .INIT_16(256'h232D3A08010100000A0C211E14303334034C4A01001F1C1D0F1F020F1309144E),
    .INIT_17(256'h48010F13071A03020806030D0505101F52610F2A203228211F2C0E11062E3116),
    .INIT_18(256'h0000000000000000000000000000000206010019607C3A1A3C682106555D0625),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_785x450_sub_000000_045 (
    .addra({addra,3'b111}),
    .clka(clka),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa(doa[53:45]));
  // address_offset=0;data_offset=54;depth=785;width=9;num_section=1;width_per_section=9;section_size=450;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hC3A6005AB3401CEAFC00CE1BF81F81804FFCC21AB098B34803800003B09E66A6),
    .INITP_01(256'hC49D1E7C42D1D7DC8A1233E235E78E03DFF8B03BAC0B0231A1E4A7F81F527E07),
    .INITP_02(256'hC7000013E0BD81FE7C649FFC80C1FCD85C07CE81803EB00803F876AC0FA7EAE7),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000009040),
    .INIT_00(256'h0400030301020401030702010502030C0701010B050301010602030700060824),
    .INIT_01(256'h0E072C25000004050300001B221443242C3940393C7A5B29111F1C0B0A0A0403),
    .INIT_02(256'h1D291C301318232933050101070342350510041C7700440C1C28032D10514B29),
    .INIT_03(256'h1C081A0C0A03120D220965442F0501001B2E305B22544C2B410F02070F110304),
    .INIT_04(256'h0F1C14070E030E2A22061905214C1F380E0001153D0C10200C190C21040F141B),
    .INIT_05(256'h1C18061E17081E1C2E1E1C181213241A342D0A2407180610385F41552406041E),
    .INIT_06(256'h28143B0A240D0C0A0324153D1C30142015090B18132F09321E1C08322B2C0F00),
    .INIT_07(256'h4B2C002B351801190B04091B071A0D001C23081F0F072200282C140D640F5134),
    .INIT_08(256'h3F30285E131E01104211310700031908100B110A090F1B1D260F0B14260F141E),
    .INIT_09(256'h180A063E362C11042A4401001C3E232302081A0D101E140508222718040E1022),
    .INIT_0A(256'h0701150C3909011037213F300205022E392B3E1715040C080A0415072C23000A),
    .INIT_0B(256'h0B07060624150A0208120C0101322D3A100601202F14522A0F042204091C0710),
    .INIT_0C(256'h37320C15120B01010D111810170F0B0B0918104C301112174B40282F471B0709),
    .INIT_0D(256'h423B090F022301030E0E0C0104070206051509111902030C67020D184308121F),
    .INIT_0E(256'h48110442335B0514141E1B101522091C111803030413262F16151A310D05091A),
    .INIT_0F(256'h183B0029431249660C41041C4637140E040F21020C210B1813251C5313100007),
    .INIT_10(256'h511400002D6729234A39081A100C1E3E2B1C0B0102041A01011005173F06030E),
    .INIT_11(256'h0116343542081441152B2E14203C02074002381505020B10130104060E0D1917),
    .INIT_12(256'h06130209071021190E0F2929023F14154B0A0E0630AE3701180806090A020207),
    .INIT_13(256'h010701200D1510042315240409012D090F08021E0E04070337163E2A000A0603),
    .INIT_14(256'h1C203433530228080E0C09091C0A0D161A2C01211D0B0400360A000851222D24),
    .INIT_15(256'h240404021A381A180F20040304220510080C0F030C1B28579B7F7D5813050001),
    .INIT_16(256'h464C1B090001000207083430220D0C060F0F1B05210001281A1C1A314D603316),
    .INIT_17(256'h26170A10090A0606040406060000171F8B455B261D0C0A03400D0C04050E0D37),
    .INIT_18(256'h0000000000000000000000000000000C0300030D202804512C20403B2D111201),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_785x450_sub_000000_054 (
    .addra({addra,3'b111}),
    .clka(clka),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa(doa[62:54]));
  // address_offset=0;data_offset=63;depth=785;width=9;num_section=1;width_per_section=9;section_size=450;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h18E0FD8F641DC8DF23CC25A3ECF21F64FFC2E037FC57FBE74F3FF7BAB290B20E),
    .INITP_01(256'hF309D0231E880021630400393870C19B06A400F076E0440E1C4140C3D00606D1),
    .INITP_02(256'h0058387003BFFF88AE3EA00D03FC40E85FE40081EC780A1FBFD0BFFFFF57DDAF),
    .INITP_03(256'h00000000000000000000000000000000000000000000000000000000000120C0),
    .INIT_00(256'h050501020801090103020201030202000501030A080602050503030005070106),
    .INIT_01(256'h000A00030706060305050129272431170F4136142A0B0C0D0400050607010201),
    .INIT_02(256'h532522084641224B3702000A011A0F41404E4B56121512115E630B202B2A392C),
    .INIT_03(256'h4721331B9F8427135B3713633D02020125264F122D060D294F1538231C403517),
    .INIT_04(256'h2B1B01072A50060705110C01121B7526320208524C0E2F071A120113080D3105),
    .INIT_05(256'h122007010008120F101D001C050C1B12230C39412B09034D551A08062007211F),
    .INIT_06(256'h162E161F04180F2B080E0D1310280C120C08000309100A4E0F48022B2339261F),
    .INIT_07(256'h3D6704054946220C05160414240D05280C212F392A090C0A1A081D2F2B5C5637),
    .INIT_08(256'h21130C0F055501250B16250C3015061239202034080F0A000B070B03060A0944),
    .INIT_09(256'h2B14041F35171F13615E07270A6928121D192433241E2A2501131533250B0320),
    .INIT_0A(256'h0E2324070F0E07071E450E1D660805620014120B080C02133819292701262B2E),
    .INIT_0B(256'h0E130E20112F260E08000C4F014F0F2A23170E5B251232091D171F12230A2949),
    .INIT_0C(256'h1010010B091D242D22120705040A2032021208563C1302062834041F2702072F),
    .INIT_0D(256'h3E1D16242713181A224B3537190C0C183926393211161F53380D060426222202),
    .INIT_0E(256'h1F0C0148092A0415161D0E04260A172F223C2C1D33290A0A2220120D1E000C1D),
    .INIT_0F(256'h35395B482D184D74332C04051102240830290112013A3C18091C11101B03420E),
    .INIT_10(256'h3F31403129431A802B3213143E207421120F0C0D40160631351603082F313928),
    .INIT_11(256'h04000D29251015322912384458270639281D4E250E0A1D175C1C2D1838072831),
    .INIT_12(256'h114312050B0C070105103A152C100008660C10213503160A2D1108110E0A1504),
    .INIT_13(256'h170A041C263E2201070E0915190C011D2F3D0639591301006E31251C10162C20),
    .INIT_14(256'h4B5F3D3C020E194B1617151A09130D12250323584637232A3705050009563321),
    .INIT_15(256'h0104090207101B59312B22703F353005080109121A25385A355A340307030B04),
    .INIT_16(256'h7D714D05000003020E05412A35361A1943490B420C3D421F243C4B0E2F988F3C),
    .INIT_17(256'h4131190D1904050100020002020202217058365749014E6D3504372C3C523A49),
    .INIT_18(256'h000000000000000000000000000000030B0003164B704D320B16323B17252937),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_785x450_sub_000000_063 (
    .addra({addra,3'b111}),
    .clka(clka),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa(doa[71:63]));
  // address_offset=0;data_offset=72;depth=785;width=9;num_section=1;width_per_section=9;section_size=450;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hE6DFAF5E10E25C40C003D609806CA0FE641E424080DC324009001803EE600FC4),
    .INITP_01(256'h0CBA191EC24541AC98F000C217866C04F003B82B633F1BF5F254BF7F3F7EFE71),
    .INITP_02(256'hC5BCD106070008677C00594A4060100CFE00C6A7A005327A0034370043EBE200),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000017CF5),
    .INIT_00(256'h0A020D010405020B0101060002030206020901040201090C0302030A05010011),
    .INIT_01(256'h1300243A070D0102010102120C0F381F30543510232C1E1E2D1C1F0909000409),
    .INIT_02(256'h0A102127546147503B03020702073550153713361D0D0A222A23063A2B816F47),
    .INIT_03(256'h00220112111B0A53622118313F040300071C4E3200292D181919000704000329),
    .INIT_04(256'h070815061D030B121619013015462E191400034A46132B3F2B0A0A0211110702),
    .INIT_05(256'h10350A150502282B300D0D1A1309030B0D0E2C0F1902054C691F160616051B0B),
    .INIT_06(256'h4210112F00080400020F0418110E2603040E0A29320232081052002E1064531F),
    .INIT_07(256'h432F12272717170716120C011C0F071E190D101C09020108070F200A353A5543),
    .INIT_08(256'h312F04380227192524132C1E191813080C1C03020C090B0204050802090C0C2C),
    .INIT_09(256'h160F210D441B18031E38016B161728184909081A06262911081308130704221E),
    .INIT_0A(256'h0A02140D102504073311020110090B6E4A3D351F091D14010517190A140F0301),
    .INIT_0B(256'h182214010A221A0B32170C13121133035B0309641616381B12040E030A042216),
    .INIT_0C(256'h070D0C1F070E0C140D0A0512190D0929111E040F481B191C280F3950310B2213),
    .INIT_0D(256'h2324090204110F0F0708040904001717000507120A0A2A2556130C0B5C160301),
    .INIT_0E(256'h1612034E1874170A17030A1405010A0D1F051B16160000081A02140B1B1C0145),
    .INIT_0F(256'h4E000E29320E13473C36431E040006001D0502191700050816053112170E3417),
    .INIT_10(256'h0F1A09150B05010C2E670A45254527191C0E2E0D171303050101180A1201151F),
    .INIT_11(256'h2F36080D0B220B0D032B281C3C3C0411480A5803000D270F231C190C210B0721),
    .INIT_12(256'h17110B14343A1D2F102A182F0B040C08601014152F62420A0E07313202001021),
    .INIT_13(256'h0A42190F10031B093750433321121523081A1963780916042D172B2118272523),
    .INIT_14(256'h041E2F468722130117220B001A1712100207380405433B8B3E0404031938002C),
    .INIT_15(256'h380808071E045D252D1228093905390401031305221A1F020B1C4A470C030603),
    .INIT_16(256'h30396015080104070C065B3A0C1E364742421B290D13040E2211231040061141),
    .INIT_17(256'h1F0620211B15000901020104020C15274C0D3016211201383D27042A070E100A),
    .INIT_18(256'h000000000000000000000000000000010003020F1631106F0551533528100E11),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_785x450_sub_000000_072 (
    .addra({addra,3'b111}),
    .clka(clka),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa(doa[80:72]));
  // address_offset=0;data_offset=81;depth=785;width=9;num_section=1;width_per_section=9;section_size=450;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hC77F004C7FE01DB0F800F118046C504000EEC72810DC1FC160E80081D414AA0B),
    .INITP_01(256'h00FBB9CC08157F63BFD1B73BFFFCE98CFD8EDFFA0BE9FF03F4FEA1F57D6F3E07),
    .INITP_02(256'hFB4430C727DC01031C1C004A014608005040032800007200BC87325FF82BCDF7),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000005B43),
    .INIT_00(256'h060C000B00060400030700010A02030A0A000102010104030106030006020302),
    .INIT_01(256'h0509170404020501040C03010B05060607070202092224081B080E0608000009),
    .INIT_02(256'h432A7D01403437181F01050403051032153C0A333B6792480F241C393B35270C),
    .INIT_03(256'h180D414E240D1021231F1E452003030B01295C270E1E041D1D1C05120216492D),
    .INIT_04(256'h333908170C04112606061A0E1A2F3F412307001F17033D3A0B0A1C42323D3D48),
    .INIT_05(256'h1A170C3E1415212A2238233A2F191B121F5206070F0606284D6539471D264A1A),
    .INIT_06(256'h272C150701131233223D10213634322B240B350B192E120C071405045411071E),
    .INIT_07(256'h150C001A0D070E06061C150E1E1D261A071F1630241D240F0A22041923100D16),
    .INIT_08(256'h260817103E110606000E1115131C200402120515190F201020182E062A131204),
    .INIT_09(256'h16192603030F081855180D2B2D294005190409132C142C1616372D1F05080610),
    .INIT_0A(256'h2C28090306001B1D190D06484000003020308186280C120B01261A1E10210512),
    .INIT_0B(256'h230F050D02040915110003081A26492C3016042B331847624B0D180C1A0E0800),
    .INIT_0C(256'h2F220A101D150318090B100114101012016E5D1A2405150E3B0F321105241A06),
    .INIT_0D(256'h62491023241D230F0F08110A100400062607010722123107190E080F6112020D),
    .INIT_0E(256'h4E0B0A0956011B2F1B000C1D16090E0C16010818111A180F0B22182450170410),
    .INIT_0F(256'h12190B0860114426542032011D0119190D17110B0C130C1D1F210A010C030C4B),
    .INIT_10(256'h1C2D0715012D0F142B240C09421839191201030211040001061A112200151911),
    .INIT_11(256'h080F0934151B0006032E4A5C4B0702021A1A3B10150A120C010311101915194D),
    .INIT_12(256'h181C0919080E1D2611351B343B145B4F61131810261A1C1A2D1F3007110F150B),
    .INIT_13(256'h1A152D16161C040A1904132922421D503209386D5F0C0408121C19160110422E),
    .INIT_14(256'h124F3647491A361016041E06120B0C3D2E2736320F1D226E42050504002F2233),
    .INIT_15(256'h1804030129093D5B310F04040F04191E06060A1C0E1C162A01140E5E01070505),
    .INIT_16(256'h11331F0700060A010303341F0E0C1F471033213916060D112D10071B1C32174F),
    .INIT_17(256'h7065200406000806020500060307235243090F13030600040C0D4A4F4D033E46),
    .INIT_18(256'h0000000000000000000000000000000605070607060041201830282619047C73),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_785x450_sub_000000_081 (
    .addra({addra,3'b111}),
    .clka(clka),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa(doa[89:81]));
  // address_offset=0;data_offset=90;depth=785;width=9;num_section=1;width_per_section=9;section_size=450;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h9877E7B01BFD8701246000BC1C01818CE00B598FBF2402FFF46EFEF8CC76F952),
    .INITP_01(256'hF28F6FFE2C227060C001000C000000C12500170A0418319C61031F80C9A37028),
    .INITP_02(256'h20730CFEF98300E2EC309C064B8164810200489E001FF7E0FDF3DFCFFF15BCFF),
    .INITP_03(256'h000000000000000000000000000000000000000000000000000000000001A13A),
    .INIT_00(256'h04020300010206030005030700040300040F09040301000C0002000901000428),
    .INIT_01(256'h0701190C0407030C0B0F02000802030005080818030607020A0C1A090A030009),
    .INIT_02(256'h1203234C6F391811040B05040003080602073D39511D520227554F3A5A5F3A29),
    .INIT_03(256'h460E03371D1E1C0F0831110D0704040704094507082417142A0B36172D280F2D),
    .INIT_04(256'h09170B1D130508000F413A1B2D86070E160808004E5C081A060E041047251C0F),
    .INIT_05(256'h0F12020F08100F0701130806071F2F161C4217040C08020810440411121F1507),
    .INIT_06(256'h0A635F2912071C23042613201F250806010F061C0B1B05031A23000637130617),
    .INIT_07(256'h011A02150D3325120F1C282B021A210C1113021B13090C071428141036250402),
    .INIT_08(256'h0203303D0817090F1E0B1F242F000C1E081114080F21141A1F0C031103245301),
    .INIT_09(256'h090B0F1F06181F121110000869254B1B043E1C0C0C18321B19302F251B0D1319),
    .INIT_0A(256'h1812100C100204200F272120081600044F223B0F1C0610191205002516012710),
    .INIT_0B(256'h151804060D1518060908222F2A4125063910080815307A13230C37000A05050E),
    .INIT_0C(256'h180A1B140412000B220212000410271021251A113F0F0E06560A19030B1B2B05),
    .INIT_0D(256'h15350A1A232C14140D020A1E350C090C161A1C190D0A1F6654010B005B382638),
    .INIT_0E(256'h2E0C10097F5308140A1A092211110B171704081F022114090D08165E220F0707),
    .INIT_0F(256'h413B0F2B210901175143161D120F0F0E03121B121F3D554C36273B0F171D2928),
    .INIT_10(256'h2E5075734D4A203F4D48000E0C2000050D062E1C070B001B0E598870729AAE78),
    .INIT_11(256'h03272705021104386A6F4253050E06190F3C26204E1B09150404222E117D5F29),
    .INIT_12(256'h320A1B040A2D1B00110E22011C29155C01040303034A360825381A051C1A0029),
    .INIT_13(256'h09090D180B12030C040D14020E041C19100B0A051E0B060001080236010F061B),
    .INIT_14(256'h471158091E1710030B0B061A0D0200040215362A1E1E30390E0000012D2B1510),
    .INIT_15(256'h1B01010409083643222E2106052514130311280B0A3A07423E33011D15010104),
    .INIT_16(256'h1F2E3F0207010A020505444D573C0810080A080A1A374014192B12341C002C00),
    .INIT_17(256'h00050109070D01010103060B0506053207190D361221111C290C321B19214107),
    .INIT_18(256'h0000000000000000000000000000000203010208354D31310D5C121B0C1A1204),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_785x450_sub_000000_090 (
    .addra({addra,3'b111}),
    .clka(clka),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa(doa[98:90]));
  // address_offset=0;data_offset=99;depth=785;width=9;num_section=1;width_per_section=9;section_size=450;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h3FF8419BFF80849FFC006CFFE4015F3F0015EF3C8612CCF1F1AF06E257196261),
    .INITP_01(256'h8B05E3BF841C7AF06F87FE22F84AC2170D0703F090F8FF022F8DF807F9DF8479),
    .INITP_02(256'h028B86101437F009B20380DC1B99FFA1C77F08BCC56A03981E2A01E3E8802434),
    .INITP_03(256'h000000000000000000000000000000000000000000000000000000000000603C),
    .INIT_00(256'h040A0A0104010409040B0208020205040A020400010206040406060200060113),
    .INIT_01(256'h0707260B020800070704080304100E0D0A01091B012A19040D04050100000306),
    .INIT_02(256'h0332322E254F221039040101000203020B1A41362B2F15154B3C48590F012635),
    .INIT_03(256'h001B140D000A28333E3D3C073A0609030F02081C401E3E291E01385516250424),
    .INIT_04(256'h2C49321C0A0A1E160C052009084A2D14380701060A1447741C216044273F240C),
    .INIT_05(256'h7C2D512C070D0B0C1B07150E080610140834042046050603372E53921D272B2D),
    .INIT_06(256'h313739615134121C0625180A12281C100B0706162F1A1A1F335F0B283B4E499E),
    .INIT_07(256'h044A011C5A64011D44402512022A1F2021060808030011171E10175627540E2F),
    .INIT_08(256'h1123144C3E260E20233F140F2D634F54041B2B390107260D071D090D1E1C1B3D),
    .INIT_09(256'h11040E002D183952430307420F1311282C4F65400847533027050705060F110B),
    .INIT_0A(256'h13020F11051503111E365F0B3612032F240F43392D193431143F480F0A060615),
    .INIT_0B(256'h233F331C0D0E0801051B091F01633832171205022231346A3C3B3B3D242A3C1E),
    .INIT_0C(256'h0F213F23013F281E0E12090A0B010F132D50191920141E1263781A0D054B8254),
    .INIT_0D(256'h861E241E2B14163F343433310B1A1F141014281D343F0E284207161581091809),
    .INIT_0E(256'h021204214145131C11030526340E0B1D17053025150913141827192913120D2E),
    .INIT_0F(256'h0A24000C07120E3531091011080700151D190F1243053D3E060B0B1D0118436A),
    .INIT_10(256'h2F06011010300C3C0E57101D3D07262640131405070402142C0C463600031206),
    .INIT_11(256'h1F0C2D0C10240514040F122D1C070413263F1813201217060B080516191E2252),
    .INIT_12(256'h07110F030F0B050A13280500080E144E1D16081A0A081904030D081506130B11),
    .INIT_13(256'h1E090B0A0013070B0B0516080B27050812161F13190B0D0401171E182A0E0601),
    .INIT_14(256'h5626051F3C000A1B081B0D060A2209050C19403A435168293B0004092F2E0A16),
    .INIT_15(256'h050006012C3F0802032C010F223A1A0405210924060E220D511607011A040400),
    .INIT_16(256'h3B66160F0011060600203B1D0E0D2C763C0B3D452A2C02340C3E6F1B05584C11),
    .INIT_17(256'h301417170F0B020008000907020105090C023F4F1B103511221C180806192616),
    .INIT_18(256'h000000000000000000000000000000060303060903083349452B2C3349021F12),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_785x450_sub_000000_099 (
    .addra({addra,3'b111}),
    .clka(clka),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa(doa[107:99]));
  // address_offset=0;data_offset=108;depth=785;width=9;num_section=1;width_per_section=9;section_size=450;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hD7003DD8780034E3E0007B14001D3EF808500F010718F2002B6519F07148298B),
    .INITP_01(256'h9CBF8119C17C86787FE2A2E7DE6D46786C1EFF8FEFFD203FFF8747FFF6682FDD),
    .INITP_02(256'h0036C761E909FDCEF8200FB0C00027B445000602802632F8C4042FEF05E3FEE3),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000005F82),
    .INIT_00(256'h07070803000F080608080B040403030A050E020206010109010F020104000102),
    .INIT_01(256'h0A050A0101020704060104000204000710404B0505120501080403090508030F),
    .INIT_02(256'h1D7140364E17351A34001108040C27330C054B650D00064A61749960242C5613),
    .INIT_03(256'h27333634151F1F2D1A0D0228310600011742393F2B3E3314071020130E3C0E04),
    .INIT_04(256'h16041142162215162232280B0528050C32090B130850501431713E221A0C1525),
    .INIT_05(256'h4D02030F4314303A47422B1A270D0C0C0703220629020508246708050A03060A),
    .INIT_06(256'h3E145563191013225D405454363828220F1D190B0010151E1A0207175A406C50),
    .INIT_07(256'h40030C0B4E1953150010252A2F2F3D3925050A150706290C1723031E2511491B),
    .INIT_08(256'h06461352101C083D74235900050A06181D070820272522410E1F04050B300438),
    .INIT_09(256'h362E3B0A2A432433496E072F603A6C0316060E2F1D160D1C31414A323030260A),
    .INIT_0A(256'h40400E01121811071E36161753110B1F1306071026222C210E032F1F383F3A13),
    .INIT_0B(256'h0508031A0D010B1003110D03121625201B1506174235070C18241D1D0B031D02),
    .INIT_0C(256'h0F120105041A1F18170825001008070214080A550C2A1100273E536519041815),
    .INIT_0D(256'h463C10150E102C251004030B000715061E04010D21070A1B0D120D0E785F5B60),
    .INIT_0E(256'h280B01290304150125083E3610041E00090F05070010120706041A510B020A1D),
    .INIT_0F(256'h110A1C013C11461E0C68313929252946380E0F030800131407000B340E12002F),
    .INIT_10(256'h140F120D031C171C4303092F2A2D23100B0516160E01010711231809390B0C0F),
    .INIT_11(256'h13061B1311010A141514041D1103062C292A0F05071A070426140B0C250B0314),
    .INIT_12(256'h01051B04050B172730121C0A041C0E271D1F0C091F140A2E090B140501110C19),
    .INIT_13(256'h100D2316021005020E0218132E1A172D31180D062C1201066D0103482109190B),
    .INIT_14(256'h170D1A014B15313D060109070E0B1D0C1A050B342A0A21423201020310176208),
    .INIT_15(256'h2302030202246B042B33211F0A100B0F030623071A0E121F1433255E040B040A),
    .INIT_16(256'h56523C0B030204050D050F180A0F04410B071F17010C0D121C0727090E403B5B),
    .INIT_17(256'h5B39110B0C0D14000404010506060500312245140D260E21292913275B435202),
    .INIT_18(256'h0000000000000000000000000000000007060603090206030C00141A19100A3D),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_785x450_sub_000000_108 (
    .addra({addra,3'b111}),
    .clka(clka),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa(doa[116:108]));
  // address_offset=0;data_offset=117;depth=785;width=9;num_section=1;width_per_section=9;section_size=450;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h71B2036C00247E4801EC06487E782661EBFFC73EE8AA0CAC0AC0290672B9944C),
    .INITP_01(256'hF14C847BDED0879FF9190D7FCD81F3FCC01F9E070F937D30E97FFF09F3DFDA3F),
    .INITP_02(256'h0754706608EF079E40F4989A8D009F98F017F8DF7DBFC06E4FF0BEE8F7D7E90B),
    .INITP_03(256'h000000000000000000000000000000000000000000000000000000000000AE04),
    .INIT_00(256'h0808050D020207070302090304060C02020F09030A03000006010107050D002E),
    .INIT_01(256'h0B0D3046010005000A0109282B2C512E1721090C11241F0D26161900050E0600),
    .INIT_02(256'h051E496C0E214D4D240208080203190D784F3D210E2600031307113B28410B22),
    .INIT_03(256'h0B0C3100303F1A505F4E6122210109011A0205612404271F18300E2231353819),
    .INIT_04(256'h0B141F0A25101102121125644010001D0002064D2C3D163E2F1610050B0F0017),
    .INIT_05(256'h011B340615030404100E16082334230012192548280F01471A15360A1A041820),
    .INIT_06(256'h0A071A0E26351F2134090D100818020E230A2E3F1E200839236B002F23094304),
    .INIT_07(256'h180C0C010F253B28023518261205010B151909031E003B1E3031192B106B492F),
    .INIT_08(256'h754F041F00260A41270C2C181C1930250F230B02021B2604152A2A37207C3D66),
    .INIT_09(256'h04170E043D0523365A4C0C092C3B062718273435041616052204121C04200F06),
    .INIT_0A(256'h082823510C08172E340E00601C0102531E6129280D0D030E13000D0B18322315),
    .INIT_0B(256'h0C0C00010E1A4725030F00046040245643001B5C436E13321C09331308020F25),
    .INIT_0C(256'h160E320F041F0E01051E2329231D081D7B22171F03070B0F52442C461E171723),
    .INIT_0D(256'hA64A2D1F2D260002110F0515060E060628070B1B2B1B2F0819010D1377161D46),
    .INIT_0E(256'h18090043A28621190E42000A0E19240B0B101F2401060B211013160C05170C1A),
    .INIT_0F(256'h160630251104205B0935012D024A0707040E2211240D16121107030216231C25),
    .INIT_10(256'h11181A0B040244140E1910263A4052104E3C1813030B00032D171A08080C0B05),
    .INIT_11(256'h010A1101103235300F0834631E4704490A32050E22354A0F1113120003142A03),
    .INIT_12(256'h0B05171B230305071307233632443332200D0E1D1A1B3917173B36120E0F1201),
    .INIT_13(256'h5C2B0D221D0F12020F0708110E0B201E3B1E3D442F070C00410F272D36050903),
    .INIT_14(256'h040805133E180B0C190F1B101F113A1203192E0C0A082D2D48010B0129273D3F),
    .INIT_15(256'h25020000090132512D0F3D380D1D1D220806062D070403001B1C1D133608040B),
    .INIT_16(256'h132E6C1D0100050306041A39151018280C2F1501220820121F020D0638160B13),
    .INIT_17(256'h10141E27260A0C020D040D0300080A361C23023228621E0226180A0F03041817),
    .INIT_18(256'h0000000000000000000000000000000004020C070A070B557B422F2C180A1129),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_785x450_sub_000000_117 (
    .addra({addra,3'b111}),
    .clka(clka),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa(doa[125:117]));
  // address_offset=0;data_offset=126;depth=785;width=9;num_section=1;width_per_section=9;section_size=450;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFCB18FE90012FE0C206FC41181B60F31F994207FC0000200B000008D8D91A4A),
    .INITP_01(256'h8F01F441D3FE023EBF202F45461EC41243EC41FE79C2FFE7BF8FFE32FC7FE36F),
    .INITP_02(256'h414767E01A1FFEECF1FE0FF165CCB9168D538921F0380A2D877680F837413F40),
    .INITP_03(256'h000000000000000000000000000000000000000000000000000000000001E404),
    .INIT_00(256'h08040607030000040501000103020104100E0D07020301000601030301060519),
    .INIT_01(256'h0F16230401000303070C061D1119422E2F56477C51674C302B110B0A03000506),
    .INIT_02(256'h280867234244271F000605000409040A482F264A28353D5546370A400C321D30),
    .INIT_03(256'h000F0E0220253B2D2316255B02060105080742335221180B030E240304082C37),
    .INIT_04(256'h260615111500032A11042736152F11650501043C191552990308050E0F010A28),
    .INIT_05(256'h21120E0A1C02170416051301001C01183148738B19040346500B687D0E150B0F),
    .INIT_06(256'h0211102C1C05151111220E030800270A151501044B5D528E2D0505260D506016),
    .INIT_07(256'h3F060210164F3F3D2B03130B20060A0229271B01060805130E4734922910070F),
    .INIT_08(256'h13496D672915003A1F48414818362E152946250824080A130C02120342454344),
    .INIT_09(256'h060502181040232A0A0500221C3B12515B2C3D5D41493B0D0D12191E00100800),
    .INIT_0A(256'h190626101B0203202E3402215D020B5F7960610D3233233D47431A141D052B20),
    .INIT_0B(256'h0F1900361003010F112028084810164260060562261E1424252B2019043B011D),
    .INIT_0C(256'h1A08111819200B0E22190412082C32100B06104A061F11250C3A3F1503090823),
    .INIT_0D(256'h23340436171A081A0001080A354E190D1115021A02012D321C120C1E33061630),
    .INIT_0E(256'h1E19000B172C0B1B030B041A09061706194A3527190304030002265205100326),
    .INIT_0F(256'h0221331926090348294E2F192D070D1519162D0918133634191C0A0531000119),
    .INIT_10(256'h201B010920091A37004C011C5A8C391108180F0215061B1905012E191D180A01),
    .INIT_11(256'h0615273E380303182B14164F2A5603150F4F23143120100E061005210E30312A),
    .INIT_12(256'h050406021306162200262231132F11041300100A1B1506243121102303010501),
    .INIT_13(256'h0E1D13021B1C170903111C1000160B15125B3B0C48080C0228321C001E3A070B),
    .INIT_14(256'h00103F000907080527281B09030721090E1914301E020D3F000001020D154D12),
    .INIT_15(256'h040204081108295A54906B31134C080022281707114F503D341338810201040A),
    .INIT_16(256'h572D00110300030501001942224A594621576B080844170F302F33150A086C57),
    .INIT_17(256'h010200000602060202050000000703060017262C19333614555F29481F002D62),
    .INIT_18(256'h0000000000000000000000000000000209070B05070C090002010002010D0007),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_785x450_sub_000000_126 (
    .addra({addra,3'b111}),
    .clka(clka),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa(doa[134:126]));
  // address_offset=0;data_offset=135;depth=785;width=9;num_section=1;width_per_section=9;section_size=450;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h1B3715E586701EFC6F1BC9CC6D3E98051BC4BDD5FFCF3B9FFFFBF7FE0A12B74A),
    .INITP_01(256'h46F033E73FE3FCE1FC1E0F24E1C091573C181D618389F2387B89030FF99831FF),
    .INITP_02(256'hF988EC9F155FC818D0F8DE06BBDFE7838EEE7940FCDECE858DC9BA6190DF81F8),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000007D33),
    .INIT_00(256'h03050501010002020001020201080600060001010B0105020102010002070412),
    .INIT_01(256'h110743490A060A07030602090F0039383332335A151C150A19081C0A0A030100),
    .INIT_02(256'h231C1843331B525C030804000A08291C18021F4B88060F521905085454495D2A),
    .INIT_03(256'h012F54140D1315071E17162600040A07271B411B45361A46731F0C011A0B0011),
    .INIT_04(256'h014B4505063701021D101D313D3E39082A010404251A1E104C252F0D11060E14),
    .INIT_05(256'h1D0101080A2A662B1306050715092151422302211C0A05134802390C181B000E),
    .INIT_06(256'h090B2E3710172325300B3B20103C15200006200D132E191A1D0D0641310A2825),
    .INIT_07(256'h14480033312A112900100B091D0864231E3618041505040A3F2114235536685E),
    .INIT_08(256'h66334432232E076559314B0F190B211A110E4B4C3426060D0D0207193A253021),
    .INIT_09(256'h08141A1D2400313A40620B05752A170A19230A201B263E5D113A14120F250D1F),
    .INIT_0A(256'h4D10312D120D0F0D1C240609570600036C3619070F0016182C372A963E052011),
    .INIT_0B(256'h0D1F1132582821230C29181811253D14090C01030D1C37142307020A22240A66),
    .INIT_0C(256'h07101E1C0823102E493C0A1B07351909323B200C1C1F05050F06071A050F2208),
    .INIT_0D(256'h593F44020F05051B0A19082321240C062C1E1B121A0D16035F0E0D001425110D),
    .INIT_0E(256'h1A0A0C176D7A222A3B011316221D0B100919270F0E0F21000F163300100E0120),
    .INIT_0F(256'h0D0B18220C054B0E3D211930040D231D2314020F040212252019031E100B0604),
    .INIT_10(256'h150A050D120B1B4F164A01483F0A5650061F251A0F051508021913122F061719),
    .INIT_11(256'h02113811111600051A1A0A221E0701234C2A3864301D120400020C0300001301),
    .INIT_12(256'h0D190D140C051729070D021F3D49104C1C120A020E4865150E0717231A01080F),
    .INIT_13(256'h371B2F21112908000503031906290E0705351E3D4F0408075E1313110B065820),
    .INIT_14(256'h1D133531631C21180F0C0705060E0B02081908132117291B0B00060658231320),
    .INIT_15(256'h1D0C040D011B130E0B175345380B1D110F090022122510160A20085A37010105),
    .INIT_16(256'h131901150902030100040027193D592010061A0024091511032128093021416A),
    .INIT_17(256'h5A010F1D2406050502050103030B02351362371E4B3415063502290F311D3832),
    .INIT_18(256'h00000000000000000000000000000009030A0207060E0C061D2058220800335C),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_785x450_sub_000000_135 (
    .addra({addra,3'b111}),
    .clka(clka),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa(doa[143:135]));
  // address_offset=0;data_offset=144;depth=785;width=9;num_section=1;width_per_section=9;section_size=450;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h86C0000B608186320FA2CB37FFCFD373FEFE3BFFFC527FFFCB1D80FC608BBF5A),
    .INITP_01(256'h7C993817EF8B68FC9CF7FF8042FFC0123FFC2363BE90460021013C0012458000),
    .INITP_02(256'h38F10010ED1D87E6CC4FC624878C61B4783A7E46007166DFB5776131D90431EE),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000014130),
    .INIT_00(256'h000507050300030206040405010606050404010106030205030504030901070A),
    .INIT_01(256'h0D0A384B02030F070200012C280B000D1D1A1D120409172C05080C0919060002),
    .INIT_02(256'h541342590A142E4D000100080711282519090D13071436334869604B2545531C),
    .INIT_03(256'h33402751502C41021B39401A020102013D350129031F18224D93834A5E3C2533),
    .INIT_04(256'h1F3D604A2949471137081104240B21581F07092D2429060605323943071E251C),
    .INIT_05(256'h232E0704100C42320313051C0E120D0A171A132B1401013E222D4340070E1216),
    .INIT_06(256'h170E29191716111A05071B08044A0D0B110F130C19310E610B3F0114492B0603),
    .INIT_07(256'h014D0C281462452A010F2D09221A30232D1B220E34093A302609180C1B663A06),
    .INIT_08(256'h373647071C2103445E0535011D09182102221C1B29424415370D2000135C5733),
    .INIT_09(256'h2E00032130101B04115201173C0B0E0B0706080A09022B12324245574A221011),
    .INIT_0A(256'h020F031A0D10171B180E1A0F570F02352E0204001B190C000D06001D284E414C),
    .INIT_0B(256'h0E1311121E10133D432E33453B07000165060C4C220F061F00151C0611151817),
    .INIT_0C(256'h0007172D1B022F172D321A0C3F3434323526060F3C050C1D1F1B052510070C0D),
    .INIT_0D(256'h0A0038070F11352001181D0301120C0628111522151D1424480A10232E04290A),
    .INIT_0E(256'h1D11086E0D1F02192219370101190B0502070B120F00100A243A2E3531160C53),
    .INIT_0F(256'h0C1022341F0B518C06202E3033182008021C0B0C110B022000061C040837151C),
    .INIT_10(256'h090F1A0F120003113C60004F5B3820040F1B0E120908070D180C0F0107090B0B),
    .INIT_11(256'h1C11090B0E052A140B060C04342F0605314B1B15061300020B140407040C0218),
    .INIT_12(256'h0A1C000C081600000210121E0C161B291609040800122B3A27092108070C0C06),
    .INIT_13(256'h200E282E0710030518080D1D111F0E002806054A0F010801520107650A293C11),
    .INIT_14(256'h0B14193A1227181B18021D0002060A2911081B173802072A2F07050303242252),
    .INIT_15(256'h270100040E1B99070008222F163A3C1B1D0E050E1A160F0A19080F03120B0202),
    .INIT_16(256'h404838030101000509042040260B09090F0E3131200B212201381B1C1A250C67),
    .INIT_17(256'h500B070F0614070902060705010B01122C175889271307041D632D100007160A),
    .INIT_18(256'h00000000000000000000000000000003070901214F42281E225B1E043E2D000E),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_785x450_sub_000000_144 (
    .addra({addra,3'b111}),
    .clka(clka),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa(doa[152:144]));
  // address_offset=0;data_offset=153;depth=785;width=9;num_section=1;width_per_section=9;section_size=450;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h970800AA781200A32044A60033BF80107FE038035C4BF03B7CC2FF06BF250904),
    .INITP_01(256'hED27FF7CE7FE7DAC5FEFC045FEF4011FFF0514F7E01A4F3CB18023C208866023),
    .INITP_02(256'h01100C00D67B018C9FA29844B81000A232001D000044C20033D19037FD1A17FF),
    .INITP_03(256'h00000000000000000000000000000000000000000000000000000000000061B0),
    .INIT_00(256'h02080409040608040B0001080002070404020006080901030109000107030340),
    .INIT_01(256'h0D030103090301010B01080305050502030A0F100405030A010500030003040A),
    .INIT_02(256'h0C2B003C303A2715010402000400050F0E121B053B537A727145242638120606),
    .INIT_03(256'h080B110F320116142558091B020001080B19182E42101046212F606F2D33161A),
    .INIT_04(256'h1008062E0E0006130A19063E1830540515080003062A0A112518061403444E36),
    .INIT_05(256'h050E0B0A0D0A030B1C060E1321052E08131E13250202040A21130342291B0104),
    .INIT_06(256'h4B121F0B0B1621162D091F02020C040B243704260B0F00531F1801060B0A1722),
    .INIT_07(256'h4E1D0B053A0414100B1313020220102C1A122316182804002A092F0602280413),
    .INIT_08(256'h00032B093E240B250A67171B18040211180C11091416121F3720041A01050226),
    .INIT_09(256'h060A1514111E2D2002090B26754C00092507020D0908233348052921082C0207),
    .INIT_0A(256'h445F110D0E271D2832031D35041604006C054C1716212F14190F181E60472122),
    .INIT_0B(256'h22104E180F36720D111A1E3025121020171A041856061A1C151E1F3A000D1D21),
    .INIT_0C(256'h2E15032B3F283002024B6F3B0510171B1D101A0723010F107240141133230643),
    .INIT_0D(256'h7D2F05123B1B1D2B28361F000C4A562202051A090C24020D00081500773B221C),
    .INIT_0E(256'h130B080D94071C1239274D2E391602120D334E450E0E11110329021D200E0A0A),
    .INIT_0F(256'h1E1331001801000E251C2A00061438131511101B10273C48001B251E20040315),
    .INIT_10(256'h09222A021223082D220306233023070D1F270217161B10301D30344C25101F13),
    .INIT_11(256'h10140A0409001501012E1A22000608242349050A20324F091A25032805301B01),
    .INIT_12(256'h0B0A122C322609282F1006011B062429050106040864050B30281C2F17290F0C),
    .INIT_13(256'h32150B081407061B0E1E0328282133253B291B01380100071B3E543C342D120E),
    .INIT_14(256'h163111141D2A1F0F1B120005070F091D26201B24320A1D351F0809050842054B),
    .INIT_15(256'h2B00000207161B483C11073B4F340F140113160205243F110C07292D05070004),
    .INIT_16(256'h1116430300010F0500151E39100B3A04062F1716040F20021D3530320B232447),
    .INIT_17(256'h3A545239311D06090005000100140121251B15580A1F08270D1B051511000621),
    .INIT_18(256'h000000000000000000000000000000000001011B511B112A3D4816043B3F5C60),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_785x450_sub_000000_153 (
    .addra({addra,3'b111}),
    .clka(clka),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa(doa[161:153]));
  // address_offset=0;data_offset=162;depth=785;width=9;num_section=1;width_per_section=9;section_size=450;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h503CAFD7914FF05EB1FE0EFA3F610FF8443ACEE0938100003A20381004641AE3),
    .INITP_01(256'h4823E146826400183E0005A3D0664A7307C1DF10F811B8FC8B7DCF81CF89E03E),
    .INITP_02(256'h06E41C680E38C017167AFE4174BBF7FE829391C2314D00327B8CA20E59C23216),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000019C4C),
    .INIT_00(256'h07010B0106070102030E06000908000001010B030A0602090301060406000405),
    .INIT_01(256'h0F07233402000A01000B012E26153F2A2411130B15210715380816020F080004),
    .INIT_02(256'h032116084A5B384B270C0101010A38062027271635683E49500C22491134333B),
    .INIT_03(256'h0C0F04407104060E583C054D260104000114081B02183D0D273D221C3E5B4C70),
    .INIT_04(256'h10070D34281B122B0E31322C61195D240702020C0902323D3A1D2C1707150F0E),
    .INIT_05(256'h1C0A050A1C201B081E476B3E344C6816431C4E2404060312464E071A2A090B1B),
    .INIT_06(256'h1D1C081B0B03031205020B131823373E626895491935701B0D220307312A1308),
    .INIT_07(256'h285F011D300A14230C000F0112170D090B23030B154F778C41021E652D1B6318),
    .INIT_08(256'h4F18071622390D37251F0F0E0801090405391A0F0B211D17291913604884121C),
    .INIT_09(256'h072A2B151B1204374970052E282F0904240A040A0B5C3C151223422020231525),
    .INIT_0A(256'h1E2B17010D04090A0D022F64300006502D000D23031F0B101242281825132C27),
    .INIT_0B(256'h100B1C1D1601312721150920240108594A040B5F3C626223053002012E16000A),
    .INIT_0C(256'h160A04080E1221170C070A06080813150E222A2E06021B1304435D0E07221D08),
    .INIT_0D(256'h3561363A13290A190A072B160C1A090814011F03041F0A0F320A190D5875582A),
    .INIT_0E(256'h1B0001333A5A060205150E0003100011210D193E1F1E1320130F091810140D1C),
    .INIT_0F(256'h171930281001214C54271A0D07250E010D141210050B1E150F121D231C09020F),
    .INIT_10(256'h260109090D06201B3951003E08272E1F130D0801000A25200C0F2A0C16050227),
    .INIT_11(256'h001D190F13051F041D1912101B260B0C10151D4C4E011608120803080A130110),
    .INIT_12(256'h1D0C030F10200D16090A0D05190D162727080607156E416B4B3303102D110204),
    .INIT_13(256'h0B150B190B140205061F040A0401161A3005321050070A046F2603271714071D),
    .INIT_14(256'h201B02254310002F120302090705091606180811180609210706020939181100),
    .INIT_15(256'h2B060305041C310F20040F262306011119170613210C0100292C4B310B050605),
    .INIT_16(256'h1D1D6D1B0C03060001013C31310446261D1F320E1200271C100222022216137F),
    .INIT_17(256'h37312C321E2B1C0B060203000014145621523B2318061E0E312C200E01032938),
    .INIT_18(256'h000000000000000000000000000000040403060542363F7627201C450B125135),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_785x450_sub_000000_162 (
    .addra({addra,3'b111}),
    .clka(clka),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa(doa[170:162]));
  // address_offset=0;data_offset=171;depth=785;width=9;num_section=1;width_per_section=9;section_size=450;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h17BC742033BF82033FF801CB06F9FEB71FF9B07FE0900A4004A000032A259425),
    .INITP_01(256'h38300F1BD500CF844219F2C456FA444F7E4A6F7781F077607987F00E10CDA160),
    .INITP_02(256'h78DB0411FC82A086A03B43E1FDA427D7FCE3FA47443F2FFE08D67D83E1033074),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000012),
    .INIT_00(256'h0004050D030902030000050407060709050203070705030001040300000B031A),
    .INIT_01(256'h18093F530808000D040102151214442E384B3D2F2C4D291B12190D0A0C000304),
    .INIT_02(256'h31171D2D2B3B4C651B030603040E30160C2A83810809121E0A400676738E884F),
    .INIT_03(256'h0E150F1D5A44455326222B2528080703190804043D2C213A1E0D3A32071F5733),
    .INIT_04(256'h140416211501110010170948281E1F3C0A0108274225160335100319001C3101),
    .INIT_05(256'h102423070D1A06130F0C1C151F03120007342C590200003023050C3104070616),
    .INIT_06(256'h22070F250009132B1004042D102A191C0C0B24232B0020493B4F0217393A053B),
    .INIT_07(256'h09620830080106022406172E44040E10001B0C220D01070619251703355D500D),
    .INIT_08(256'h0220022D293B0A3F670C13080A081411090807181E0B092107100115013F2C0C),
    .INIT_09(256'h0C07070B260D021709240B252711360C0D12131D030914222B2F0A0421141115),
    .INIT_0A(256'h0B0B4147180E12053702241B3210094E012A24131417030A1505110E343F2648),
    .INIT_0B(256'h17121B2D253D0C162E07081605090E035B041F330C243D430512200A32061B25),
    .INIT_0C(256'h3B0B0B0200040100091D181303040D01060C02493B020E181910400E050B0B23),
    .INIT_0D(256'h161F32053C2709031D340E030C0210080A193C171F1A2F4D04031508216C1238),
    .INIT_0E(256'h1C0C0B0430071B022F260D113E2C220B07060F081C181206111F032401190D1E),
    .INIT_0F(256'h100E0B3D1201562E472D022813301307504C331F011B17150B0C110E0604220B),
    .INIT_10(256'h2627200000053258485F005E6B27222B001A1D113C31382B241F371B06081306),
    .INIT_11(256'h27211506010616372F0616332D330127300D3715170E01220F0A19463A140723),
    .INIT_12(256'h05090E001702110A1906071539020D32201604011D203505161A1A06120A0B17),
    .INIT_13(256'h1110043311080C19100D020C1814151C1F1F123E0203020668190F191911271B),
    .INIT_14(256'h0D4A19041A0500584103030C120F14282B0C0A1F2B281E3714020401382B1234),
    .INIT_15(256'h19000206242A631C06060820212C1E050F0300161A120A020F160A2A210C0502),
    .INIT_16(256'h1A26040403040000030E5F29170B2D02070D15130B031018140D0A0310131104),
    .INIT_17(256'h3A0220170B1A060B06020003010E202D310C4C9607023329154A15121531201B),
    .INIT_18(256'h00000000000000000000000000000000010000154E6C450D346E1A0D2922030F),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_785x450_sub_000000_171 (
    .addra({addra,3'b111}),
    .clka(clka),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa(doa[179:171]));
  // address_offset=0;data_offset=180;depth=785;width=9;num_section=1;width_per_section=9;section_size=450;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h60AF1F7F7181FF721A5FE520FFEE30F37BE43781E456C7AF241076EA444AB208),
    .INITP_01(256'hDE506781C01E2F27BF830057FC30B4BF84AE93A406E50BC8EF587E1DF706E8F7),
    .INITP_02(256'h3DA93842C1F8E1FF2EAFDC58784C078EC01E7C388CBDC02087BA02837CCCF938),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000001400),
    .INIT_00(256'h0005050204040300000802000806080008020A030A0405000804050104030328),
    .INIT_01(256'h13040B0507010900050004030A0A0F0F00393C1A0B0C02050201040303000303),
    .INIT_02(256'h34261355052533381D0501010002130E01033F613E241B180F1D301C08321701),
    .INIT_03(256'h021E2E3B7D0B0A554A4D172700020205170D251B091C504F04140D100A070519),
    .INIT_04(256'h250A220A0C131C4E74390F0E14080A4005000D420F2F08561A0E1D21230D0D1F),
    .INIT_05(256'h020A36080201020300220D236FA6200C32AC20291F180334262131071514421C),
    .INIT_06(256'h8F3D4D0605150E061C01020E0F1C440C484E18371E3D4E46046D0C1547110E05),
    .INIT_07(256'h005404342518313D06000A29010A031A0B312C1D6547310335165F591F642802),
    .INIT_08(256'h5603631B250B023415512E182B02060812260A130627120D20244927161D915C),
    .INIT_09(256'h060D2D00482A341F580200560E451504000A282B1E09051F12111D0416080028),
    .INIT_0A(256'h1C00062E0C0B0416151C1F014B01080A602636351D0736201824231804080404),
    .INIT_0B(256'h100D1F18110A15051508100A031E250B0B041E0A381450621101140217080E0F),
    .INIT_0C(256'h4E5B523015031A1320141413080C081B0B0D52211E041402071E84A265604D27),
    .INIT_0D(256'h491C0C34132B030D28090D0C241E060707070D220A3111154A030F061D0B3B54),
    .INIT_0E(256'h1D100204004A0B1D581602131E1C09201E0C0C00150C0F0B132C141F04190509),
    .INIT_0F(256'h1B073B070C0C0B021B2200162800230D0C1F1C182D0B0F1F1408170B20291D12),
    .INIT_10(256'h0E0B1E343911122F5B55092B011A2F130D131211240C0A0C1D0F0C1B14111514),
    .INIT_11(256'h1D15100914110C3D0D05023731010134163F5E181D1B160312162A0C0A0A050C),
    .INIT_12(256'h0A27160A13011A1514030D19091523602701150D3849522D05300217082B2D0F),
    .INIT_13(256'h7F103F34081E1E030D0403080F030D1319252E79550709092616102D5617072F),
    .INIT_14(256'h05555C1A333D342D050715040D230F00140E152427121D171E0601070A182D2A),
    .INIT_15(256'h0009010B08060E0B1E5310120145020E181E0F01180515030920062811060104),
    .INIT_16(256'h4758491E06020902070B483E1D262E1113160116160F0A08100B352C358A4A2E),
    .INIT_17(256'h4C382522090200060A0004070100000B1D3A26302C31251D081D282825241016),
    .INIT_18(256'h00000000000000000000000000000001000105030205040F5030306B6A435348),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_785x450_sub_000000_180 (
    .addra({addra,3'b111}),
    .clka(clka),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa(doa[188:180]));
  // address_offset=0;data_offset=189;depth=785;width=9;num_section=1;width_per_section=9;section_size=450;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h800098F20005AB31443C170687B86012E7E910E7E0A8002E03A00000290809C9),
    .INITP_01(256'hABE07C0E9D4FF3FBD80C2F9D80C151FE04E627F7C1627FF83487FF814C07F00D),
    .INITP_02(256'h79207CA707C388019CF00200BF6000162C07C98040782C02F0438C3D943C85FD),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000006FF8),
    .INIT_00(256'h0601010208070106010006070104030108020B06040402090408070A03090111),
    .INIT_01(256'h0C042011000102030200010D09132C382E455A81715F51161D1D131313020300),
    .INIT_02(256'h26483840136312150D03050301011942232A2E5A5C714D240A000F2F39592345),
    .INIT_03(256'h221B0915120A4958413C27361C0005062C1B1A100D5B693B0E011B0E0319481A),
    .INIT_04(256'h1508141B0C0505050C0C0905140A0C281D030502142E12221437110311070504),
    .INIT_05(256'h071B05212604091B12060A2403120A07062F1B17450201203537232B02171D02),
    .INIT_06(256'h242524190D0C223B2F2727170D0B120801040214061E211F3910010149822D06),
    .INIT_07(256'h5F030E044D0F2527221C1C1A102826090707190B0A0E030D290249112C00050C),
    .INIT_08(256'h1A07290E2D05012A373111082B2420381E25290A04241407020418000B03191D),
    .INIT_09(256'h16080D250B0631181B08022E7314508047654676695F542C1E161B0C2423000D),
    .INIT_0A(256'h150E0E240C0610190007190912060806407A7DCB876F7B4E4A573722131C0A14),
    .INIT_0B(256'h01100316081E010C0B050C100612300B0B000809086CA75C5960411B0B16101E),
    .INIT_0C(256'h190427090506202801350B150A0F1A04054E0012091D1710174F13245632040C),
    .INIT_0D(256'h622C2F0C0D1B2807291503060932001D110602140F100D44181613166E441108),
    .INIT_0E(256'h30070D352B0D301E0E0A152B1C0A0C0A060704011421022C2C0C204C111F0C20),
    .INIT_0F(256'h200105442D0905602C41060D2A2F41270B11101E240B0409111619032E0D432A),
    .INIT_10(256'h13010211010A21524316076C4904141406264815030406131F01071D090B0110),
    .INIT_11(256'h1C0A352216441C00000C0F3B1B0E08308D086D2613052C061021011836020315),
    .INIT_12(256'h04051C1504050F0D0208180917002421150501034F1546311B101D22300B1000),
    .INIT_13(256'h0813042301090D1C1109222202131603250C24023B07060A0209210911143628),
    .INIT_14(256'h1B120102131D0A0222010112181615240D02042A1B33263B1403000116080A24),
    .INIT_15(256'h0808000618332A060B20381D0D1C1C181411130E241304280B063C5A18020405),
    .INIT_16(256'h2E5F640E0704030307096038363511041F1D1C241654632E49814A3A244B3620),
    .INIT_17(256'h120E231F1B060105040703040903021B1411604C887323180F22021F1556621C),
    .INIT_18(256'h0000000000000000000000000000000000050500241530473D1F3F3005100026),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_785x450_sub_000000_189 (
    .addra({addra,3'b111}),
    .clka(clka),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa(doa[197:189]));
  // address_offset=0;data_offset=198;depth=785;width=9;num_section=1;width_per_section=9;section_size=450;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFE1F82DCB3FC58EE3FF708E07F6C67C14013BEC826698C00090402E31012F8EC),
    .INITP_01(256'hAE8000FC40A004641E90CA40E80A2C062190993B1A4F8E36B1BE814737F85FDA),
    .INITP_02(256'hFF57FFFF1B4FFFFF81FFFFF071F1504666A10024422E060006C623026FC8201B),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000010FFF),
    .INIT_00(256'h070807060A0E00000300070D02030E0003061106090204020805020607060108),
    .INIT_01(256'h13031B41010001030701051C200106130E1C384B030A07060C02030A11070705),
    .INIT_02(256'h01511043381D3D2F320407080303260709081D131531265A2F1F114C605B5C33),
    .INIT_03(256'h0D0400073D4C3C266B612B5A3000080C16031B0A05134800200E1326011F0F28),
    .INIT_04(256'h00090E2421180909201B060403222E0C2609052A07555F382236073505131019),
    .INIT_05(256'h1B040F180633312D250C070E00102825120C3E1F2F19022A214C011C1B361213),
    .INIT_06(256'h5F171D0A12290627081A372F0706200A04110602110C63082D4E062A3B1C2120),
    .INIT_07(256'h2F6D07112B5B4D0F0B2C180D1B082C300B0021060414100B250106163F3E5D2B),
    .INIT_08(256'h0440042C0B0C1653425839221A2814090A040C1D070505060A0F01040F120602),
    .INIT_09(256'h1C040409041F200D4D6004261A6E040B1B0B000B08180A0E140E020B04051120),
    .INIT_0A(256'h063C1A19021113011C0B00156D13014B340F270D0508041C0F100106140E1000),
    .INIT_0B(256'h0C001509061F1B0320250E0A2D0200275B041E544C2585031E05060812060D20),
    .INIT_0C(256'h0B311A080306040D191E300706150B062B1A183C15151618110C35191C1F1B05),
    .INIT_0D(256'h0A3E2A10183A11160D0A20092733270311090A00060A42513F0A0B1775362C10),
    .INIT_0E(256'h3D0E005027603A1A0C00230F030B17052B0B04200B0205320308094D2C050333),
    .INIT_0F(256'h0B000C0A0201427830161C1C314111241F030C052B1121131626020605070D15),
    .INIT_10(256'h15051A01140D1C0D575E0D7324711D1D171301002815000B1520250D0F02090A),
    .INIT_11(256'h071820170C0A04250D08001539410445785A2E1A170D011815221424201E0405),
    .INIT_12(256'h0B0708191F08040A220015021A430643590F100C5312320D0F37300C1E2A1D15),
    .INIT_13(256'h1A080B211E08100B090C18010510030B0F28162D5F030C00730B1734230D2012),
    .INIT_14(256'h3330290F2515001A09110A19100A0C150203161B0404000C400300093A32161F),
    .INIT_15(256'h070903001B490D1E1809314559502055182E36283925322B1E412302180D0004),
    .INIT_16(256'h19241E1803000A0B041024242B639FBC9C613C4799761C58665A2F443B0D0455),
    .INIT_17(256'h792B131320110A0200020D0201031C0B838D8F69500D1583594B4D45347F9048),
    .INIT_18(256'h00000000000000000000000000000003090000003924232E56544F47624E607D),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_785x450_sub_000000_198 (
    .addra({addra,3'b111}),
    .clka(clka),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa(doa[206:198]));
  // address_offset=0;data_offset=207;depth=785;width=9;num_section=1;width_per_section=9;section_size=450;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h19DA601119C902D7FC0C0E7B0364BF843FDA60236009692006400800E06F91A8),
    .INITP_01(256'h159D86195A8CE91DB21C04DD31E015F0DE0D360CE050B00E010184E8100FEE05),
    .INITP_02(256'h002F00328881C780EDD8F313ECC7D0A1E0329B1387B1ABF6799199A711199A71),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000008010),
    .INIT_00(256'h05060107080605000306010A0301080103010905040000060500030402060520),
    .INIT_01(256'h140F302D09050200070B0C17131E312920300438062D24223816240C06060B00),
    .INIT_02(256'h09112852561C435404010207060317090317131202220601516A0C1D24323646),
    .INIT_03(256'h192606211A0F160401250B011905090009153A560147213D290012081C650C04),
    .INIT_04(256'h0D1211071813040E0C0704151B0A1710160102010C777B172517201817041921),
    .INIT_05(256'h1E27011C1E150A050F030A0C250E1F120E29252104050A00016E644127172429),
    .INIT_06(256'h062807230F06140A0D0A170008010902080B12140E2E120B0D1C05070B111B56),
    .INIT_07(256'h0A120213443F1E23350D0034230904080A20040F020C001F1F0902152126490C),
    .INIT_08(256'h0D1F3D2D2607001F090030011E260835181801020A24141420120F1809080704),
    .INIT_09(256'h0D22101E33300B284C6800041650300308021401020426191A2D221A081F0A1D),
    .INIT_0A(256'h19462423191E2128090D0F1B3C1D010B180B05050F4A240A191D2814062D3410),
    .INIT_0B(256'h0A0B0D0322262C013E2406160F051B17290E02032F071B012C39100006012002),
    .INIT_0C(256'h14230603200D1E145426052530372024112B0F344202152750201B040C152500),
    .INIT_0D(256'h111F0108041509002116141E4D2E0033122E13390403210C06140C020F020E19),
    .INIT_0E(256'h1710034D51220E031E0A0901170A29262D4F2B20012A320A060D1E3E20090D2C),
    .INIT_0F(256'h00231A0E0704065603051028080C142204052C2910665F08171E1B2803220320),
    .INIT_10(256'h162F070C1B053214176101392A030C1F12191832020019243D385C1F02190525),
    .INIT_11(256'h0412372B0D1C1501021D2E1818180011264103231419000201060232283B4409),
    .INIT_12(256'h0D06192219112417090104050225191041110100244433321C071D0A19050918),
    .INIT_13(256'h28050602051518241604100D060505031E2220255402080160510F0F09191822),
    .INIT_14(256'h200220020A010E0311050F10120A03391903102217193E1B3C0405092529011B),
    .INIT_15(256'h340701050F30300B220F1002090810052106113103122A2E1B6A431300010902),
    .INIT_16(256'h020838030900000006006C7C5B4600110A0C020C1A22293C56271E2E31120315),
    .INIT_17(256'h442229171A0C0404070205000601254E1B2031481A0B06180B023610052A1F41),
    .INIT_18(256'h000000000000000000000000000000030303001C3B685D0D195B010F14200348),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_785x450_sub_000000_207 (
    .addra({addra,3'b111}),
    .clka(clka),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa(doa[215:207]));
  // address_offset=0;data_offset=216;depth=785;width=9;num_section=1;width_per_section=9;section_size=450;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hE03F0A9F628519D0C0513981056E1800008743CD3D67C1BFF81FF77FF4E10D7E),
    .INITP_01(256'h07E1040552B003E73F800C5BF80FE87C00E699C01E0F1EC591F48E45BD2A40B7),
    .INITP_02(256'hCEF2FFEF1F4000330201006D000E187001EFCBA062844204314F00C700CC9C03),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000011EFF),
    .INIT_00(256'h030D0108030101050104070600010103080001010406000C02020E0305010B21),
    .INIT_01(256'h0F11425104040002060B001A291A39331E423A3B1E403A13051815110A0F0406),
    .INIT_02(256'h0F1311381231054B1B070F0402114137111F00210E28281D1F1613523A271454),
    .INIT_03(256'h2F1E2529300B1A1C1B11091F27050307080A08342209021511040B1D32290905),
    .INIT_04(256'h0225300F1B060A080E1226160C330C4F070204492933431D324A180531173D40),
    .INIT_05(256'h0F26040C1222121309140710052305011311113F0401083E2E34002132331808),
    .INIT_06(256'h6B322C000C00030E0E0811070606031609051509094B254F254B0C2640010A3C),
    .INIT_07(256'h1D57061A2F2C0209070D06060B06070B01190A050A0C23050C2A29093556691E),
    .INIT_08(256'h061C012C390D01450E3F3309021C0D0A0D0E0E050604090B0515020D0A050A2C),
    .INIT_09(256'h21050E05201211181771033B44030508130611150203130B04013A030C081410),
    .INIT_0A(256'h183625101F1C0A0C0F0B07212F0E0B4BBA4702171602141B0606100E10082028),
    .INIT_0B(256'h0C281629252937131E17120B0A0213126301205B1D12040E1D130D1903110F20),
    .INIT_0C(256'h14170C0A082F2A162B1C1804020E06080301060044011217030624091423110E),
    .INIT_0D(256'h301F3D0B1B251308110F2B0F22181C19230F0B0610022000480A11031B43161C),
    .INIT_0E(256'h2C0A021A0A492305120C07050A190E09130719201D15041B131912223D05101A),
    .INIT_0F(256'h210F1E1F150E44231A090506132C0F04020B150601011621212B1F0002060402),
    .INIT_10(256'h271316040D100041596B050D41023F1D10132506201A13161B06001404250413),
    .INIT_11(256'h15001B110B2424110E100F0F2756040B0B4627340D2225070B1D0E1312024A0D),
    .INIT_12(256'h0E021D19110618081A2E2012110D05172C0C080D151502513C3D572600081717),
    .INIT_13(256'h4350312425030008030511031D171111201E091D170502047420063C474B5F24),
    .INIT_14(256'h513B2F432356262B221C100003060C000B1A2D0317061A554206020A000E2432),
    .INIT_15(256'h2100080500321A231A2F2F2A3900100E14011329123123130E531A3711060001),
    .INIT_16(256'h213C380C0108010105084A6B31292103220C1A350A2503010D04050614040751),
    .INIT_17(256'h5715070E0E08070006020305050008076D3A43702E17020E1E3D122014232922),
    .INIT_18(256'h000000000000000000000000000000080806091654594004467816044A3A0D31),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_785x450_sub_000000_216 (
    .addra({addra,3'b111}),
    .clka(clka),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa(doa[224:216]));
  // address_offset=0;data_offset=225;depth=785;width=9;num_section=1;width_per_section=9;section_size=450;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h87FFFFFABFE02F09FE00307833C1A7BB391A720302AF00000960080106018C96),
    .INITP_01(256'h89FDE3523F543031F34086341400A40041B040002D80801398A8A7EDDA47FFDD),
    .INITP_02(256'h6178009FF27C7DF097FDFD14FDDF91B7DB9218F840C5CB9C1E8787814033FA1F),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000004385),
    .INIT_00(256'h05070200050A07010200020602050001030B1108040A0501030301040001010C),
    .INIT_01(256'h181E23180100040806040B213027524627452176012B5246431F131A12050404),
    .INIT_02(256'h0D1E52873D1F15022B0002020B020C1C161218373239594F383A0E812A3D605F),
    .INIT_03(256'h23032E260B002706284248372D0303000A0B280B080A0C3C31071C5700231D17),
    .INIT_04(256'h211E021006100A070B052742483543661A0907220C77783E0D190D03130A1107),
    .INIT_05(256'h4A61310A1C0F07180612162C0D182B2C0412091B0904031E59072D1F1E0D232F),
    .INIT_06(256'h2F330A52734853352A28110809010D0C1E14211B211B23430E2104140C7D0F21),
    .INIT_07(256'h286C0019471E3C2A44222C20482E3A32411A1F0C0A15280202230E414C11060D),
    .INIT_08(256'h111B0E2606440446050D08000F103A2B202B394F341E27042B260002321F220A),
    .INIT_09(256'h0A011216120C43151F17024C2405403822280800010D04101017180923081106),
    .INIT_0A(256'h4213150006040709011B32322202005921362D1019141B094120120B21012E07),
    .INIT_0B(256'h170A0316181D11141D0612230022214F6A0B0E642E4219200A2101083C372D14),
    .INIT_0C(256'h232D150B0516110A242920090416050019061A5F3B0A002D1F2E4F2E19000F2F),
    .INIT_0D(256'h40081821072503020602272544450710130B1212070C4832260406021417001A),
    .INIT_0E(256'h060F035325100C01010209010A070F194427170E000002091B0E0B034015020C),
    .INIT_0F(256'h041E0D26120F0076010F04240B160C0C0504080B1D121D0D0A0524042723221C),
    .INIT_10(256'h010F0509060D34073B330310365B16130A01031913250805070D093E10201104),
    .INIT_11(256'h252C0912121303100206471C0A1D011B533B0B021410030D1D1C291D1F0E0008),
    .INIT_12(256'h1801070F2F37220E0915172435121D054D01050B3521150A282829011417101D),
    .INIT_13(256'h5014150F09241414180503120E0102250C101B126C030A00240A336C2A1C4629),
    .INIT_14(256'h0A2773710413230A20161216263539553F1E060D290F65264707070300378E81),
    .INIT_15(256'h0F050D031D0C636B2F24314E3425090120171C4F370B15242021204510010603),
    .INIT_16(256'h1D271C070E040203071422334944041D1B0C21424C3B1B1D58272214091A3C32),
    .INIT_17(256'h290802000408160203040703050404462A0B4E3E302C1D30023B0D06305A4016),
    .INIT_18(256'h00000000000000000000000000000001030602051D2324204334452228100B02),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_785x450_sub_000000_225 (
    .addra({addra,3'b111}),
    .clka(clka),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa(doa[233:225]));
  // address_offset=0;data_offset=234;depth=785;width=9;num_section=1;width_per_section=9;section_size=450;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h7F21FC16A01F68CF01392AC00F912B407911A787EE030FC6890790E0D1A77451),
    .INITP_01(256'hE01E096905D1BA91703B976700F81E602FE59607FB50A01F9F7B01F9A1F01F80),
    .INITP_02(256'h036C0E30072DD618485EC2134EEC47ED0FC038921C1800A1C001BE0C0E8DA0EA),
    .INITP_03(256'h00000000000000000000000000000000000000000000000000000000000170FC),
    .INIT_00(256'h0401000301020001020406000401030500050401020606000002000605000309),
    .INIT_01(256'h0405352F0500030507060010140A1E0F0714250710051C081C0E110507060401),
    .INIT_02(256'h2252401709105900090508000601103622225A63110206010F27158C49242013),
    .INIT_03(256'h0D10081F142225171D2E3E4021000302054A150725112A46171F0D071E21320C),
    .INIT_04(256'h1314050007081C1201162B0928251B0F0005013D33002C0E271416000D35300B),
    .INIT_05(256'h113215041D28021E040E082207060C0A000526733909014010040D281B0F1D2E),
    .INIT_06(256'hA303090A19170B352134092B15050D210A031406031C3348063C002959305522),
    .INIT_07(256'h260D0601A0053E06210B0D2F3A322A123526212011041B061212150556193D23),
    .INIT_08(256'h06030F0C0E0E0803752211111902143A314440195D3020320B01131F29023114),
    .INIT_09(256'h041204160E01312C5D490A0954072C0A320E1C2E20463B14442C251D280A0302),
    .INIT_0A(256'h21150B220B0014242001103C120300004503170423193B2118030503452A1210),
    .INIT_0B(256'h15001B040110192B070D021A2E062D2E1800000D345517292606101E040C1D11),
    .INIT_0C(256'h2521373E2A2B0109030E121B2A12072A070634360D0C0C002F693B1620050927),
    .INIT_0D(256'h580C0A13051016252314010313030D2D10133801071405222C0B0C055F382002),
    .INIT_0E(256'h1614002234090C161C141C021C230909200D031D2106040E0802085938140102),
    .INIT_0F(256'h150F1C122314104017170F28302016051A071A1B0D0203140318180D0C040803),
    .INIT_10(256'h0B15080002251C120D3C0C04201A0F371506120428251B2001060C000715040A),
    .INIT_11(256'h092913291200000815072B430D3605021416180D0804051A0A2319142C14190A),
    .INIT_12(256'h130016130C0C0E171D0600010805074A36321615064A18050B1302200F17130F),
    .INIT_13(256'h140C0B090203040E0A1101220600060D0521191A15061305480E1B010F080F06),
    .INIT_14(256'h06062B030216061007281017280F0716100E041017174734320106060A131C10),
    .INIT_15(256'h0D0A000302252A42260C0C1A222935030C211A0D110B02120037296003000506),
    .INIT_16(256'h35265A150B060105002823020317210D3B4117240F131A222E43210B235A6211),
    .INIT_17(256'h432F212716000702000B0A0706082E3D8C61040209241900160312074C200642),
    .INIT_18(256'h0000000000000000000000000000000E02070813334838242935470F1A5F2336),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_785x450_sub_000000_234 (
    .addra({addra,3'b111}),
    .clka(clka),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa(doa[242:234]));
  // address_offset=0;data_offset=243;depth=785;width=9;num_section=1;width_per_section=9;section_size=450;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h6F7401F7FC809F2D9807F82C38FC5661FEC4FFFFDE51FFFFF41FFFFD29AFE352),
    .INITP_01(256'hF17FE1CF3FFE01F37F8009BFC211FA7031F3F2073F1F00D3C0F01C7C0F008405),
    .INITP_02(256'h06E4100009BC00012E07B00685F20739576E03BB4F6138067F95A47FFF533FEF),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000013E60),
    .INIT_00(256'h0102020905070007020402030604070202090A00050905030102000408000305),
    .INIT_01(256'h16050601050B010105020233290F0C110F130C0B070A040F1206141A18020006),
    .INIT_02(256'h653A3D0E3A370C0A0A0406010304021E26112A2A2E0856604E707A642326463E),
    .INIT_03(256'h392A272C587F030E103D4340130408040D102F3161691C318E72694497873F5D),
    .INIT_04(256'h0C00262B22031D14393D480D262B150A0C060001212D163C221E07282D040037),
    .INIT_05(256'h35070F09060F160C18380D17100C120C40692B110801020A46320C03010A2E13),
    .INIT_06(256'h3658106E460B120D0D05091B293B360502001816113B3936311704060E020230),
    .INIT_07(256'h0D1806095F132D2F001402071A1205080B171D0C000F20170F0C19044E230117),
    .INIT_08(256'h28111A3E390F06190B1F061016031506070B0E050001181F16211D0426030702),
    .INIT_09(256'h0B0A13320E131104033207442938305E52001C100D1F0D000F10021D0D0D2420),
    .INIT_0A(256'h150F2B2816150903142B280403020B0945434367612319030802020F0F05061A),
    .INIT_0B(256'h05020D1C00300E18130F19040F16012E49150C092D0715473E3C310C03090E10),
    .INIT_0C(256'h2B09160309120A03003010010C1904031016050335151012190F1911182F2A0E),
    .INIT_0D(256'h0CC84A450A171826010F03171E1F372835372B0023060834160B0D1004642E2C),
    .INIT_0E(256'h1313042F598C0B3108082019111D07201E3D391524100A172F1E05640F270706),
    .INIT_0F(256'h1C43143B5115322815012D26270827250F222E070E452D1211170B0C442B2B16),
    .INIT_10(256'h1E53663439110C274521001F360593040E0B020608032D110301041708282217),
    .INIT_11(256'h1E0D2D3C342A22160C0C150E400B012D03156807200600131808130306122A55),
    .INIT_12(256'h1902071A0528070906252D17251523105309090121700B2A2C02050009060407),
    .INIT_13(256'h010C0D22021E1E040A1C0F00010C122D2A10291834000F082931051C040F0404),
    .INIT_14(256'h292A2E2A160D0D1A18322A0D06081A120200293406010E0F42000101203F120C),
    .INIT_15(256'h370101000E2B233B33371916082350100A0F0B011E06152D210C6B2F0C040C05),
    .INIT_16(256'h333A3F1E02040E04050746392C122036120A1B0D27410214421D2828084F1E63),
    .INIT_17(256'h00072428191F190408020109040F2E472631220444522D2356242F40411B1C47),
    .INIT_18(256'h0000000000000000000000000000000503030801070F1C29194137061A072421),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_785x450_sub_000000_243 (
    .addra({addra,3'b111}),
    .clka(clka),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa(doa[251:243]));
  // address_offset=0;data_offset=252;depth=785;width=9;num_section=1;width_per_section=9;section_size=450;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h1B305EC44FB5AE046E0020CFB760EC2EFFBCBDFE6FAF0FFC3059201F1E52181D),
    .INITP_01(256'hFB6E00BDBFC00BF9F901CF9F8B01A0F9007E0730058A7291D803083CC0D897C7),
    .INITP_02(256'hF9F8BFFF36CEFFC892CF3C211FF009977EC70177FFC0C7F83E0A3F25B817F809),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000007BFF),
    .INIT_00(256'h000D0302010C0B020B01010402000600000C1203030203000006070103050012),
    .INIT_01(256'h0F00171C030404070006010203161701090E281C365227000512050301070801),
    .INIT_02(256'h049C74363A132A3D0D03010307134F431310000617085E3122252D03353A211C),
    .INIT_03(256'h130629072E4C6E15230E02020B0206001E150A2A2146032C2B1E3A1A1E431007),
    .INIT_04(256'h100604050F1A11270D0439203137002A040201432709153432170417101A0902),
    .INIT_05(256'h03061100130E10010C18160A2916030A181234241808014913044D2512283C11),
    .INIT_06(256'h6A4225370F161F14040A0A1210070912010D230F330438665C29031E1922720C),
    .INIT_07(256'h3D55061115180A4208100D1700141303010D08050403261A1F1611777F1E6424),
    .INIT_08(256'h0E1F1A02404B072B2315070502071E20101B240A081615021D040C180B03224B),
    .INIT_09(256'h24392105132B3335246A020E203C160823032E1E060C0C0419111C0A3B270819),
    .INIT_0A(256'h2645531A042F120B3C1E15110903024551355C09130002000617080615190F0D),
    .INIT_0B(256'h020B0510172A2B241C0404171602080D0E0300490505592100090C1B010B1823),
    .INIT_0C(256'h12400100050E100D102941160A272934210B23202A1C00032F2345453E1C0B0E),
    .INIT_0D(256'h4B2B3B2D2208180B1B27070A1D11330A15030C0731220B55260A030886023E47),
    .INIT_0E(256'h5125023F60732D1E483E1A0B1E15210B2039240A14030C3429050753361D001E),
    .INIT_0F(256'h3B1303492C2351721C3F4C00483E070A16291B0A1D1E141307140E1B4213045B),
    .INIT_10(256'h240504020F252C10024A0C2E45263C494D2124400F031304122E1A0E0C00062E),
    .INIT_11(256'h0F0812011B040B0100184713254F011215390F3B54191A4D020E02071B04090F),
    .INIT_12(256'h240D121301041C141008110F27150A35150807132954568305282D39050E0202),
    .INIT_13(256'h47268A372A1E190E10020807100603090B0A060E090011036B11013D1A39354B),
    .INIT_14(256'h412C14500C16555549251C07141A0717000E1A2610060C390807070175282F4A),
    .INIT_15(256'h05030406212A4B0101021D0B50513217100C16180D0F02120D46083430000208),
    .INIT_16(256'h181B18160A06010308083F3C0603120F2A5A593C52321C0C2907040013332867),
    .INIT_17(256'h1217322B1527120205020407030B100207030A40684A2F27806F40383D300E02),
    .INIT_18(256'h00000000000000000000000000000005000902020507021148352D659638490C),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_785x450_sub_000000_252 (
    .addra({addra,3'b111}),
    .clka(clka),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa(doa[260:252]));
  // address_offset=0;data_offset=261;depth=785;width=9;num_section=1;width_per_section=9;section_size=450;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h20504261842E631400FC153407A0D100CAEC291278BCF7FFC87F81F97632F052),
    .INITP_01(256'h1E499E21EC0AD41F807F81DC13181D203B00B0038007033046907E030101B07E),
    .INITP_02(256'hC685EF8FC5C3FE7E3FFC1D82BF1058237800067FA006FFF30199D92432347866),
    .INITP_03(256'h000000000000000000000000000000000000000000000000000000000001BEFD),
    .INIT_00(256'h05090207000701000701080407080A0F0A0206010506030500030001090A0617),
    .INIT_01(256'h0C103B40010300050402021B24082D2214232B060A1608082605140B09020305),
    .INIT_02(256'h0019307A291760452F00050803021639263A434E1B2C7D87978859609C875A27),
    .INIT_03(256'h190C100010181F181C1F2C0E2F0D06051E15060B11302628001D13262B190601),
    .INIT_04(256'h0812060F18081101200C01154E350D2F1C0602283C3820031916081D0C030C20),
    .INIT_05(256'h2A0F241E1E1412150C04050311241E0A5D8C430739160128333E174606080B11),
    .INIT_06(256'h09314A60100301262B19010A2B1B2610031502113C421B1E260008300F13041F),
    .INIT_07(256'h5832073A17165925270A17150D0F231A021B0D04140C14082C1913415010691F),
    .INIT_08(256'h070106214202041134585C1004030C19211011160E0B0D0D1C061211112F4A10),
    .INIT_09(256'h0008061012120F460768023821050916400B211E100609001C060E031F160306),
    .INIT_0A(256'h0A080404000C13261B0A28630D02033F823F39120F000A080813161518150E0D),
    .INIT_0B(256'h210C170F10000521001D2D301C02575A3B090943271002200F09032708121F08),
    .INIT_0C(256'h0D1F01091B03340B0111020B091B3227202A1C223408071F10240A0C1A0A0110),
    .INIT_0D(256'h86004920171B17061E042D0617161927080A16231D39196C11050F1E6703050A),
    .INIT_0E(256'h2B0E052F971902020A103A070A1104002127003600152D1C1116311C1E0F011D),
    .INIT_0F(256'h0916151D0E110F611D02091F040E2C0121251D0C13120C000418151008203A05),
    .INIT_10(256'h0F0608140E1C0711193C051F0024151B030E05040201211700140329180B1201),
    .INIT_11(256'h0F36181B280A0E1008160D090F4C080E115800330804030D1E1E02010B031901),
    .INIT_12(256'h1F100C140020020902060E0D000803163C15141110703A300F150709070E100A),
    .INIT_13(256'h142927050E00000A161A280D101F0E072A0407281B1013076915451C031A2923),
    .INIT_14(256'h26302D0C31393B320B0F0A10110F1A1A1316140B121E0705100607024F031D2D),
    .INIT_15(256'h0C040C0122511422315A296919251400173C0818220B070B24192B3C0604020B),
    .INIT_16(256'h471B3002000701010D0B533E130B27425D201626690C251E1D3E562A2C6E361B),
    .INIT_17(256'h1B0A091A090B03010D0301030306010451701B202E43827813283E3F2623013F),
    .INIT_18(256'h000000000000000000000000000000060204080B4262401945530B112D171403),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_785x450_sub_000000_261 (
    .addra({addra,3'b111}),
    .clka(clka),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa(doa[269:261]));
  // address_offset=0;data_offset=270;depth=785;width=9;num_section=1;width_per_section=9;section_size=450;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hC5827134D8045E42C10DD7A4C20182760F0FFB09D52A003311023F82C22FCF45),
    .INITP_01(256'hC5BF2FFF3DF007F26DB03F1D741131F9C013C7D613F44F136F41FF80EF77F331),
    .INITP_02(256'h480E010220B331E383BBD20C6202304E99401DFD0001C9706085A057F87B0F7F),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000005FE2),
    .INIT_00(256'h030100080302030004040E020A0603080B0B020B0404070A00080C0104010608),
    .INIT_01(256'h0000090C07000205050806000504050005030C0B040B06060503020000000509),
    .INIT_02(256'h3B2D0A0913040F0D0005050B0305085758567557605B4F482839322208080B04),
    .INIT_03(256'h24200A221B182215111D1E2E1A0304020415152C39050C330000030A0327171F),
    .INIT_04(256'h1B1D0D11090703171A00050A1E2C1F341A0304002E2916161301160823240D2D),
    .INIT_05(256'h0A06040A0200030D1419071F0326260D23200C09410D0D280A2A1C070D281102),
    .INIT_06(256'h01013E18040324351E0F15012102051811170F0E0F212F173912062C14120905),
    .INIT_07(256'h5006040A0042001E010C0E08270F08101706070E040000101F1F25062A070846),
    .INIT_08(256'h23101E253B040D030A100421280A192B274950170F00090400140A091D081301),
    .INIT_09(256'h08080115240A0837240A0209353621201A170B322C224918020010070E02210A),
    .INIT_0A(256'h0D2E130E010A060A261120590309053945100B03201D070B0C1D0C0F1A19081A),
    .INIT_0B(256'h0F0F07011F0636211B0B0309131B163D0905191E333F13122811120C1C180B00),
    .INIT_0C(256'h0024110C061504001B0926021212100B261B1249011713124556082217000B09),
    .INIT_0D(256'h3B31041C020D0006100D0A1016193008270D1E1C0B2B2711112012137D621406),
    .INIT_0E(256'h1C28020862250914250B130721010904021D34300C2F785C5643224B06110400),
    .INIT_0F(256'h302E1A29380A3906372A0526201C1C1F17000D07061033388A8272495359492B),
    .INIT_10(256'h3F040621140032464E5C021F6F2E45200A250002011E021801466B806B48284C),
    .INIT_11(256'h1807030401100E05240A27241F0605296F550F00141C0B0C071600050B174240),
    .INIT_12(256'h07080C0D08093C28050C463E092F570F3C1C0F035B2D32240C091A0A010A0808),
    .INIT_13(256'h320F260B01040A09060220221A06250E284A3D08560600054E0B0C2C29021F0E),
    .INIT_14(256'h294A341F1705080D121A060B200402122D0E080D21425C442805040615152718),
    .INIT_15(256'h030102072626482E1D410A151304331C130708041E210C291A21155D0A030409),
    .INIT_16(256'h5A2C2115030600010A1916083100012D030C130224581E04091839094A311909),
    .INIT_17(256'h00170602090D01010E050005010103324B2E42292E212721184E010E02181033),
    .INIT_18(256'h0000000000000000000000000000000B0A0B040530362708070803155E422F0E),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_785x450_sub_000000_270 (
    .addra({addra,3'b111}),
    .clka(clka),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa(doa[278:270]));
  // address_offset=0;data_offset=279;depth=785;width=9;num_section=1;width_per_section=9;section_size=450;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h90FC368F9F83643DFC2EC7FF81C00FEE8502CFCCE4381E152A0767FCC2E48227),
    .INITP_01(256'h9BC25B8E9525C0634218963E0D7962E870251E0F02E9E1E06E823E1F288F83A2),
    .INITP_02(256'h7999E60FF1E0F6C0131F7224FF6C3C8F76F481765DBE0C67C22F867C29DE1593),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000009BDF),
    .INIT_00(256'h050400020002030007090103050A030503060001020603010302040B0102040A),
    .INIT_01(256'h1000070F03040904030900170B011B0A1D1A180D38233A26020B030201010205),
    .INIT_02(256'h284E0A622B041B2C3700090C030408255E4B0E11354C140E1D5C1A13180C0A25),
    .INIT_03(256'h0A1D0A04001B162203337457380607013513503D032943254B1A1C0B151E0619),
    .INIT_04(256'h170713412E24151411100C0A0500273C1900020D4314334D5D241D08310E0B00),
    .INIT_05(256'h1C46592F22180B20121704091D0D030C0802454C390502045235113A2E184E2D),
    .INIT_06(256'h141D0910377F333D1500142F2A09030C041725200204495416280239312E0E24),
    .INIT_07(256'h8C07040D21122809519D5F171A102258280A2523000627073800213742010140),
    .INIT_08(256'h08183B324C0A0F15103708401759AC4B1F0320794A0E202C200410111C2E2203),
    .INIT_09(256'h00060A0137060B4648130059250A2E2440083A6171200B3A6639040E10153A02),
    .INIT_0A(256'h29230B03061C020C301804063C08002717194B0A25240942615344194B2F2E1A),
    .INIT_0B(256'h0102071F0F0D0215132409071A0A0303140715468F34471718100504395D4912),
    .INIT_0C(256'h091E0B2D090602220A03181E09161A250F2E362801031927935E4D0117002229),
    .INIT_0D(256'h4020040F2709041003020530010612170A2A0F27160B54511805191008171201),
    .INIT_0E(256'h550C052B0B122A0410081D0000150615180E054221420B370608365900150A0F),
    .INIT_0F(256'h1F03141A65200258010C0E0330380D0700100D1201230B110625120D173C1208),
    .INIT_10(256'h28270401141B1218462B0C09400E1A04290D060107031B0A2543121009171034),
    .INIT_11(256'h02112012212A18212700130333550A081827070B0D2115001D1E0B13090F0A02),
    .INIT_12(256'h1C010305191E090B08050207031C1C145C0E04020E352109071010003E030318),
    .INIT_13(256'h0A0E16071A1F170B0F0D03030C02082C0802465749100402052538100C2D2909),
    .INIT_14(256'h0543487A05341302080B22092014130E051817070B0351471A07060602385435),
    .INIT_15(256'h010201012930010427390010310E250C15310709072B101D0F2F092915040000),
    .INIT_16(256'h404B4B0A040C000B01022222130F2207114B41010558182B4A1D081B44110E06),
    .INIT_17(256'h03141B1712030406020500080205021F5F7513374504143D11090D2824532A50),
    .INIT_18(256'h000000000000000000000000000000000400010A0309061C312803044D192712),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_785x450_sub_000000_279 (
    .addra({addra,3'b111}),
    .clka(clka),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa(doa[287:279]));
  // address_offset=0;data_offset=288;depth=785;width=9;num_section=1;width_per_section=9;section_size=450;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hE8F8CFF51F98F371784FA60130FEA0877FD812FF8CC8BFD13CFF9C5E611F7E2A),
    .INITP_01(256'h0EBB0003428084040E1C0040FD860C03B14C157F0FC3FBF97431BB0F871D68FC),
    .INITP_02(256'h86B3FFFE110FFFF94DFDF0F44E7C1225CFC24725BF081340E0160007004B6040),
    .INITP_03(256'h000000000000000000000000000000000000000000000000000000000000CDF8),
    .INIT_00(256'h010101080603060300000005040303030906090C03010300090101070202040A),
    .INIT_01(256'h010F0309010F05000409010F181B3C2507222C4A0F1009270602000508040102),
    .INIT_02(256'h2026250B04084B09160300020405284A1A02243C041C3B34203F340322362429),
    .INIT_03(256'h0E213743260929142113260727040006290107150B2D101203010A262E060312),
    .INIT_04(256'h1809071516070D13324141370A25202C15000828243C3E140B27190706071E06),
    .INIT_05(256'h0B140E05030A0906100B190D224C272118074811461303244523101D180D1C0A),
    .INIT_06(256'h361417042E0B210C0E1D08010214092A23522B110B172A4C545D032D2B371606),
    .INIT_07(256'h170F0209072B3300282113061B0B0E00080230301D3C45290A1D053F082A5527),
    .INIT_08(256'h042E1319210E0C25020C3124141404240A0909030C161C130837501547273541),
    .INIT_09(256'h0119260426080420166807540F1E15231D0E04321C0422080715392403163A1D),
    .INIT_0A(256'h0B0412030D150715231818224B19042E083B152A09071406180E2A30151C250C),
    .INIT_0B(256'h0F030D01031024011120070D26170D3D0C1209353A0A0D1A1A051404130F273A),
    .INIT_0C(256'h030612030E0103191E082F0307030318110013480B1315144F001D14210F0F13),
    .INIT_0D(256'h195A47140B060915051710112E0A2A0A0014000F0B061D5303100F236B313825),
    .INIT_0E(256'h2A16055F768D0601012C14181C3E1012030321230206110C061004240021033E),
    .INIT_0F(256'h2B0A1416031C5393052B2532020612131C1B26250F0B04130112280D21080D09),
    .INIT_10(256'h0002191A13000829275F016A121A061700060E120C06292A16170703000C1C24),
    .INIT_11(256'h1B07180A002749120A21030E450505464B0706222E1A1A18281426301404210E),
    .INIT_12(256'h160A1002110D040D10362C12171E1104271E04023A20050207131029150F0606),
    .INIT_13(256'h091603320904040B300A140E1D2C0208010B003F3F0401046727230D2F190D0C),
    .INIT_14(256'h261F031A0E282804082A2F09161514052D1300231904213E0B000B025C380E05),
    .INIT_15(256'h0708000A0A1B3D345E2409090352010B261E18010323151318332F0D06010C06),
    .INIT_16(256'h4B625315000400010B093E2A424C77401A455142835F510C6E659C522E223A18),
    .INIT_17(256'h1E0F1914001307040402010500000E4C3406144E411C24807A0E2305622E351B),
    .INIT_18(256'h00000000000000000000000000000008040402010604160A0D03090B24033801),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_785x450_sub_000000_288 (
    .addra({addra,3'b111}),
    .clka(clka),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa(doa[296:288]));
  // address_offset=0;data_offset=297;depth=785;width=9;num_section=1;width_per_section=9;section_size=450;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h8015E19447FE1B607FC1B68B9E1D00DB01DE03F8F399200838A8760D4CEA1234),
    .INITP_01(256'h4F1773DDFBF81F9CE3E2049E2020B880483FB10081F903CC159401E1DC001E1D),
    .INITP_02(256'hF92ABBBF134200708C1D03F2E39416857DC0EE47F01FFFE707E98FB0DEE0F71D),
    .INITP_03(256'h00000000000000000000000000000000000000000000000000000000000080FB),
    .INIT_00(256'h000200011004050203080B0203010704091113070504040B050002080502001B),
    .INIT_01(256'h0F1035430101090109000408030C2D172421272D340C0C04401D11000C020106),
    .INIT_02(256'h0311161F030B3B4E13000408070808170D140638746C434E99512F06172A2E22),
    .INIT_03(256'h0619433920091A0947352206090405000D2A5F41001A84847F70260609173635),
    .INIT_04(256'h06250035224310133427320509400D10000700451E5B3A450A0A011C01051828),
    .INIT_05(256'h05163409282221072626092109380C3220171C502209024901370A1B2D132016),
    .INIT_06(256'h4E0F0F21170716300F151B0F20220C0F404B1926430625433B1E082700372124),
    .INIT_07(256'h312C0A1752431F2301040D220504011D203F1B1E262A0408100E1912582C2733),
    .INIT_08(256'h271332010A0F0111034C1322132318210A0400151F3D19281E191B2438101B30),
    .INIT_09(256'h1E491B1C0829051301500310050949101025050705080902322B152C30340B0D),
    .INIT_0A(256'h200E331E1604040913453A19320C0E622B1C231A16111A1518061303161C2729),
    .INIT_0B(256'h1A0111021904141420080E1104145A2A4E0A0B54013247021F0B0515060D0B0C),
    .INIT_0C(256'h493F111C130825180C060702180E0D060419351A0906111A081C141C302C372E),
    .INIT_0D(256'h02133507001C11050112072A2B0307090708041D0007020B3F0E0C0A47080D21),
    .INIT_0E(256'h4B0104273A2021131C21451E1203020C0E0D08180A13062009000F144D050208),
    .INIT_0F(256'h0E1729305106531040621F03070814070F030A0E081D090D2829001F14183309),
    .INIT_10(256'h09030A2933320A34433913165B475307072D28111B052F18221C292A2219200E),
    .INIT_11(256'h0A2F283F0A0514035752792B2504031B03144B19052036190D01461130151814),
    .INIT_12(256'h061B110A0E040F2700102C023F45761A290B0B20272D21431420080003212401),
    .INIT_13(256'h01061E08181E0C0B141814201F1D22172A4C54081A0F0A022B0D1D110A02060E),
    .INIT_14(256'h14280E3965380C28250010070C08060A252D140A01610E13020502070C200203),
    .INIT_15(256'h2A0004000F1C1A2D551100042E091E17060F102210140C180A3D54042B020701),
    .INIT_16(256'h0C2D0623030002030717284A443E06022B1C0A5823210C1C0717241C16003026),
    .INIT_17(256'h060C1F291A2C10010002010504041208301130340300343B1E21132B430E1E44),
    .INIT_18(256'h0000000000000000000000000000000404000615130A0800331A252B2205241F),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_785x450_sub_000000_297 (
    .addra({addra,3'b111}),
    .clka(clka),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa(doa[305:297]));
  // address_offset=0;data_offset=306;depth=785;width=9;num_section=1;width_per_section=9;section_size=450;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h56600340B609F5E3E4E7EBB10176BF4E0A59E1823EB0FC01C41FC0A423F1220B),
    .INITP_01(256'h1C3FF60763AA60749248126218C43C650017341F9A7901E3CF86063CCF40F37C),
    .INITP_02(256'hF8A01FF7C23FFE07C3FF003FFDFC038D47F025637F00260EF00062FF052073F0),
    .INITP_03(256'h00000000000000000000000000000000000000000000000000000000000190C3),
    .INIT_00(256'h060104010004060306070D01020001050B06040008010C080400010A0101040C),
    .INIT_01(256'h1402423C06050002000001020B10150605033440093413021403020502060000),
    .INIT_02(256'h221B4319161E353B06070403000A342F0F20181C6645083C6389924E151B1502),
    .INIT_03(256'h1C15191703090412391F3434050505063D09133A4947061401081E0D422D0619),
    .INIT_04(256'h0F150D181E1A0B030E092910410910090D010B4935410C2E09191D1B11180906),
    .INIT_05(256'h012E140B0E010A0D080209060B1D16240A3E28582803013D1E08022C080F0B03),
    .INIT_06(256'h10241D131F010319010B0800100C00060127350901145339241F021116063E27),
    .INIT_07(256'h41120045122B2910020C02160E2202000700051A0F0C2904161702123F20090E),
    .INIT_08(256'h0520161320160908070A1B1D2529391E180B120808150901160314070F4B021E),
    .INIT_09(256'h29280049142E32195159042E1A5010182A32070A1310270F11050E0E0D110D23),
    .INIT_0A(256'h101E0C040100241908565A185202001B1D1D26391D0E160A1627260C3118141F),
    .INIT_0B(256'h07060A07042421210D030D1F1045473E0016023008132D34391A021F35020816),
    .INIT_0C(256'h031900190806150008050F25190E080D0E172C38131B000A6203111F19050C1A),
    .INIT_0D(256'h530A0E2C0321130D0D18200012000606211B0E08071845141718050348051C0A),
    .INIT_0E(256'h18200167220F2C2911201800130519050413053145514030051B3B340714072B),
    .INIT_0F(256'h2C150C0F1816007F16121D190B060B09131615150A0B1516465735161E020323),
    .INIT_10(256'h00653A1B1C09130D163007466C27121F020B0D100C011322113958221959371D),
    .INIT_11(256'h3625304D00232F2D0A0B0A0D434701146914261A1E1C130A140404061D23606F),
    .INIT_12(256'h060618251C0E3526102B13343405174F401507074A554833190B081618282501),
    .INIT_13(256'h0405071E050E2F3420100A12190F13253533181A440102010F44073632111502),
    .INIT_14(256'h1F541E38292402042E402C181E1C090B0801280F050F0D2447030700114E0D31),
    .INIT_15(256'h06040B000E373E4B456C4B634D243F2B04191E050919303E4505463D100D0401),
    .INIT_16(256'h2322000104080D030B0F4A405A52464A41351C122A0D1A295A50504F5351341E),
    .INIT_17(256'h152D38391C090A070A0B01020A0015132100174367631E0E0D2B3E23180D130D),
    .INIT_18(256'h000000000000000000000000000000030100000D3F615C35010E392F39302A1A),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_785x450_sub_000000_306 (
    .addra({addra,3'b111}),
    .clka(clka),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa(doa[314:306]));
  // address_offset=0;data_offset=315;depth=785;width=9;num_section=1;width_per_section=9;section_size=450;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h8701FD98900798A883F1C8487F3C26408E2E88004284014404700C0282190B13),
    .INITP_01(256'hA8EA1FE88D47E0934475993C0A092343A0C1DE70267703067F7C7C67C341CF70),
    .INITP_02(256'h060D830CC47CFF0307FFD10C9FE89863FE08E01C000F898003BBBE01E317F8FE),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000004E00),
    .INIT_00(256'h02000204060805020006070109000001030A010407060A0C010104050505010F),
    .INIT_01(256'h07044B490E050606030101020A22422C0E361F3407151205060E180A11060900),
    .INIT_02(256'h1C2526310243044815040B000004231D331627320E23371107070B2D200B0228),
    .INIT_03(256'h120D1E17020B07081E54010A0E060203070B3D110E0C3A2E3439313C1C0E220D),
    .INIT_04(256'h060D13130D202A0B1103264944261C5E1C01024C452C1134002804101A2E150D),
    .INIT_05(256'h292231030F130C2D210733230C2E1C382E1E425D4510004643141E0614184A3A),
    .INIT_06(256'h0C1A480501123921151F1A160B1B2635400C1D181F12431E6314012E1F205E18),
    .INIT_07(256'h5123041B60340F0A332D2C0B00271D0B05031F1E2931091B16473E0F580E3935),
    .INIT_08(256'h340D11081E3507350920261B2505120816010E0A0F1117120432140F043F5205),
    .INIT_09(256'h292825064A241D012A0304402B3B114A4506053A141D111E2316030D280F3823),
    .INIT_0A(256'h40101B180B0C160E05060F11270C054F231C180B2A0117221110082038073A1E),
    .INIT_0B(256'h0D0403152B09190C0E0212072707070C1204165022192224360410250D200D18),
    .INIT_0C(256'h0723140B0B000203200812020327001302130910090E03080013112B22111A02),
    .INIT_0D(256'h059D040C32021201041507270201370E0C1415040120054143180C161E55170C),
    .INIT_0E(256'h231B00074F7C2422221020081A2B0F282A2F0F001B290A07071404021D210622),
    .INIT_0F(256'h09011C000718553802BA5503100F040D0D1900171F2E412215170C251C030117),
    .INIT_10(256'h041E110A171E200F185E03180664540D0705251B1212281806324719180E0310),
    .INIT_11(256'h392435112528010603140A02265208251C2F29010113070C1C1B1E130E0F1802),
    .INIT_12(256'h0E062A1E36272E111110140D123F3A0206030B0913263943120000020F19060D),
    .INIT_13(256'h565C6936311F111B241E1F190530140A050C0A16030B0309020C2B458F370027),
    .INIT_14(256'h072E346327448C5C313E3E07140A04190613180A3415001D4F010C09011B4019),
    .INIT_15(256'h2300000006271B291D1B3A99753A462D5034040C0D020609161D5D3C090A0404),
    .INIT_16(256'h0A230A1403040C0103035A6139200F071206134C45462C1E02323F1A3A0B2B3E),
    .INIT_17(256'h01041923083124030002120105170044321A060D08082C0A350C0014010A0124),
    .INIT_18(256'h0000000000000000000000000000000402060204010304033E3619316E25190A),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_785x450_sub_000000_315 (
    .addra({addra,3'b111}),
    .clka(clka),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa(doa[323:315]));
  // address_offset=0;data_offset=324;depth=785;width=9;num_section=1;width_per_section=9;section_size=450;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h1641F7885C04E004263821C31C4F170004F29C059BAFF013F20FFFFD90D0E7F8),
    .INITP_01(256'h02F00620258048026800800028080003E81B217207F0BF63FF83A0FFE1001FFE),
    .INITP_02(256'hFFC7FFF3F57F2CF8E3970CC67FEA282F2CCF82FC9FF637F1FFED7D0FB86F91B9),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000018F1B),
    .INIT_00(256'h01000A01010400030104000203060003020A0A020101010303060503010D000D),
    .INIT_01(256'h1307464201030109040101000924442C1C361D74013B5B2921101905050B0109),
    .INIT_02(256'h281A02554408644C0503020101172A4E190103183B767530121E2A0F3C36363C),
    .INIT_03(256'h15082C211C0720072C4B43191500040404340F7732020D14333744421E16191B),
    .INIT_04(256'h22031D1B14041528061C29231C385D3D0C010A04076A426B24251D242E160E0F),
    .INIT_05(256'h001906170E1A020D0800021E2502172B4238021A0E0907080F0B06090D011A01),
    .INIT_06(256'h0B64101D0A20100000030B0615070E101C3007243357426B2E2905333A240201),
    .INIT_07(256'h3C100008200F191A10191D0118070C01212A350B111645171C152B621617023A),
    .INIT_08(256'h3724381D7D10014A3E2603061712040B0D1013262036273C1F20123B42080E54),
    .INIT_09(256'h0D2B1417293A49521A0A001C4953072A1101170A0C091C0E133438443E392A34),
    .INIT_0A(256'h142219123B0C110C25095225040A08031902170F032E280D0710010D29042717),
    .INIT_0B(256'h0B0C01020A13212829191907050C26123D01051F12270C211422221800000D01),
    .INIT_0C(256'h0F091805190212001F0D1F08012C2A1C3C370C11350B082425333807131A0615),
    .INIT_0D(256'h4F0E020C082B181F191823261A1F2411020A12394E46227F3115091F2C101A1D),
    .INIT_0E(256'h4A11072962042E111F5715382F3A172F1F090107052C23432D3933864C170234),
    .INIT_0F(256'h0E281A354A202B191B0D1C04185015082317141A060223020F1F060D1C274448),
    .INIT_10(256'h160A101D1B001223143008432329050203341B0D150D1D060A14201E0B1C0F0E),
    .INIT_11(256'h3918251F25322101152918371C4601242F2A141C12040B260000090320142E19),
    .INIT_12(256'h070601101D3D180E0930050D090E2A4F571F02082E01141323181129030C0718),
    .INIT_13(256'h0605071D261B000614100000022F180B0D0D3A6157010C0017466214010F0B0D),
    .INIT_14(256'h104B46352D07401A231F20040503010516040443091E3D5B4700020311484D0C),
    .INIT_15(256'h0A0101020C116B6F4B0D150A0205091A1609171403011A1E172C2B202E050B05),
    .INIT_16(256'h7848310C0504050702023E1637270E28060C0213030E171C1C55272E1E043100),
    .INIT_17(256'h46362F3A26030706020504000607242D12265B4D08160C0A0A20191519050787),
    .INIT_18(256'h00000000000000000000000000000003020001020A040B0E555D0E3F4410644C),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_785x450_sub_000000_324 (
    .addra({addra,3'b111}),
    .clka(clka),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa(doa[332:324]));
  // address_offset=0;data_offset=333;depth=785;width=9;num_section=1;width_per_section=9;section_size=450;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h01700E660C8027248226737C05E6348E00E05C000C6640BFC930CDE84FC4FD2B),
    .INITP_01(256'h18FF0FC19FD0F609FD0FE107F03FE1FF87FE53E07FC90E03ED50112649032186),
    .INITP_02(256'h42127C007ACEC00B6FFC9FE79FFBFF1BFA4FF9EF29E7CFF170389E07011FD070),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000E12),
    .INIT_00(256'h061201130101070204020004050504050B0B07040109010E01010104060E0108),
    .INIT_01(256'h15160C09060100010100050804101E16210D016B0E37071113010A0204080005),
    .INIT_02(256'h5339640E6B51543A320802000006440A16151F34101F3907112F0C11113D241B),
    .INIT_03(256'h1640200702112E145A6E394C3A0700020911340F5220550E32381F1E01153B24),
    .INIT_04(256'h03350A110015000D242B323A0C397E3B1D00030D39163D054E05060A01130B13),
    .INIT_05(256'h15011C22161007000A021403010B30011A1A3E2310060708134F1D1920171112),
    .INIT_06(256'h8A241C292134070F031413231D062F03170A121320414B311225040C59121F0F),
    .INIT_07(256'h302314534D5F4B05000D08100916041D1928290C02211F2C081953074B0A512B),
    .INIT_08(256'h07580B0F222C082C2F95231E2B081C2500210A1C301A0607042103150A1E1F03),
    .INIT_09(256'h1136390A02441F08214907382443392F1B0612030F170609132A030C00152A01),
    .INIT_0A(256'h2D134E1E11091E04382E4D2A120E09095121040120170E042B3712221B12241D),
    .INIT_0B(256'h12220C0B250F39162E1D032E2421121E060A01090700593636120F042E17033F),
    .INIT_0C(256'h96030203000F070A1A0D1D0C232E18292606202C1C161F091A46848676071D15),
    .INIT_0D(256'h2E437D41552C180A24050E070F0E093A292C150510402619081011001B194F48),
    .INIT_0E(256'h40290211133D197444551306091704070902253601050B051526531627180407),
    .INIT_0F(256'h041B0B3A171144120B771342765810041D310E1501071B33260D01310B1A2107),
    .INIT_10(256'h031E273C2025013E0968121116250C3A5F1A0B08082C16211A192D080A061D2B),
    .INIT_11(256'h0318192302000B071B010D1F373A010D2E05321E36292013222409000D0E0D05),
    .INIT_12(256'h21110D0B21080506161A1A0F0B1D1F1220100C1A30AC0C0D1B264C0625240402),
    .INIT_13(256'h75676D2F0D110100021303090E2C1207022C2D103B090507610541095B3F5313),
    .INIT_14(256'h230D38636F5E16281C120606130334072139130D452113162F0A03094911467A),
    .INIT_15(256'h05030B0006332F37A3992152781508171F01170112191D173E2D363224020205),
    .INIT_16(256'h032A38080200010202051D4D1833183719151D10174140101A6264311B003412),
    .INIT_17(256'h32062B281F10020003020209030109324707102D2C0921221753263F636A884C),
    .INIT_18(256'h00000000000000000000000000000001000905020F020C010F3130114A2A0E46),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_785x450_sub_000000_333 (
    .addra({addra,3'b111}),
    .clka(clka),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa(doa[341:333]));
  // address_offset=0;data_offset=342;depth=785;width=9;num_section=1;width_per_section=9;section_size=450;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h178301803DF99482BB98C808FD8061EFC00706B3C0022F0005C0200092708423),
    .INITP_01(256'hC35E106C3DE402C104407C3AE00FC3E200D40F003F2AF807F8AFA0FCA0B91800),
    .INITP_02(256'hF8A177FC787FB3D9D384EF058029BF12067C3976D34E065E7EC0BDC1ED138387),
    .INITP_03(256'h000000000000000000000000000000000000000000000000000000000000CF11),
    .INIT_00(256'h010B0305030104090B0404090B000200080E0202040304050106020400050507),
    .INIT_01(256'h07000707030501010401032728203219121A0E372A17160017100D0402000000),
    .INIT_02(256'h180A5A73001308081E000006030116023C452300053649412A71214F1C425E3E),
    .INIT_03(256'h351E10122214571516524749390105041800032C03210D160401053621143F49),
    .INIT_04(256'h053D370C060406051303222A0338213420060A4345230F172927201924060D46),
    .INIT_05(256'h39181A2321011111190D0D0F0E1C041D0340202E2C10033D19325E1621000214),
    .INIT_06(256'h150F0616301600160C0B1A0307101A0F0F0B010F0A1956352045013115311B05),
    .INIT_07(256'h854904103D0B284922100B0A050706280323200022231D020A175F465B175B2D),
    .INIT_08(256'h03000F7F2E220E290A14371D4E141401184D29090C030E0A200B1C1605061564),
    .INIT_09(256'h061C0D0814320B9B0967045C081F59461F04022224352E050C0D230401020510),
    .INIT_0A(256'h0A1C072015181C0A003D0B59050305422C2B965E0D134D201A14160D02101C16),
    .INIT_0B(256'h2C30303E0E0702002C13081B01110E363C0D082B4E4D582D1D0F0C10132C3E27),
    .INIT_0C(256'h18011011001C12091219210B02092828401402433816091B2A083410372A1A0A),
    .INIT_0D(256'h2A211405061912250107221E3C2D16230C05255347310C3C560B0F16474F0A18),
    .INIT_0E(256'h0A1C023D0A29281D1704210B0E0C0D05301A0C4014040C020D4A173C21220A15),
    .INIT_0F(256'h26180019581D166E3726040D1F0C19060212001E2813160F102109093D414724),
    .INIT_10(256'h02070105240A261F55590827281228370802090D1008080D11360002001D0809),
    .INIT_11(256'h242607060D2905073417450B0139011919100D0D0A0F0909130F030C0A1D0410),
    .INIT_12(256'h0D1805060801101305120A030A1F063718060002093111000503060B08160801),
    .INIT_13(256'h332E11080F0F052700040D12110215050815211406090F034D09322013031400),
    .INIT_14(256'h12531B0C0A1C23282C140415010D0B0A0E040E143A243B402703000329390508),
    .INIT_15(256'h0D030C011F142E0A0F07161C0A100107120F13101427201F353D091228070107),
    .INIT_16(256'h1308421302090000080744423E5E211D0905062C00001237100F142E1F4A3B17),
    .INIT_17(256'h0D151A1B0D1906070800040407010C1523013B2F19053A492A3B292A0321070F),
    .INIT_18(256'h0000000000000000000000000000000605080C09091B0B111E4E020102221007),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_785x450_sub_000000_342 (
    .addra({addra,3'b111}),
    .clka(clka),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa(doa[350:342]));
  // address_offset=0;data_offset=351;depth=785;width=9;num_section=1;width_per_section=9;section_size=450;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h464AFE48707FECA6E7FFCBC20F8037808073A048362B05EF749F06CA88425007),
    .INITP_01(256'hF08C107F65BD0FE45FF0FE443F3F447D77B001E77872F86600A02300402B2700),
    .INITP_02(256'h008ADFFEEB7CA1C68100177E000059006208800C405403C000041E000505C007),
    .INITP_03(256'h000000000000000000000000000000000000000000000000000000000000FDC2),
    .INIT_00(256'h040305010D02020B0206050600090400030204050D0A0106080B03090201021F),
    .INIT_01(256'h040F0E0306060505040005020F101804000E1E151E0E0B000D08060103000602),
    .INIT_02(256'h368603242D2C181C2B0108000303070E04353E2F0A15241742373C030F12221F),
    .INIT_03(256'h12000017316C4E24022534203A00010F0304192D322D0C312322000C20171C38),
    .INIT_04(256'h0B00250F0E1E1D3D280B14211316663A2901013917090B01010B282C09222804),
    .INIT_05(256'h03060E130018101C0B0C14152641471325281C404A0A013B0B05040721201605),
    .INIT_06(256'h22132504200C09160801030F17151D46073D20122F2122143C4C031D0904111E),
    .INIT_07(256'h1D2505345541251C0D061B2010000C040C16152621191B3314071D0D5F594A2E),
    .INIT_08(256'h26191521381B0722BA1C324008000309000908100C080A0707030F1C10083400),
    .INIT_09(256'h19071C483A141E3B032E025962161120192503030E02200308070A3534051915),
    .INIT_0A(256'h163829301D22134D1C0705073C090C5701180F15010A10150608210A05132810),
    .INIT_0B(256'h0E051F0C12193E342C050F060207041651011657312708260C09060C050C131B),
    .INIT_0C(256'h0307241E200A1D150E270B485744313300212334350A001B2D2A28341F2D000A),
    .INIT_0D(256'h084C260E061B4141131B072C1838390742646326140D0F03180E020A2E051917),
    .INIT_0E(256'h1A04041C12100F020C024B0411101E150A302E201A2D3D2B4D3E391632100B24),
    .INIT_0F(256'h24110A200F06032609021A370F03112E0C0D1B05263438420F14354940330B08),
    .INIT_10(256'h0D05100D101110032313003C0F0706343A3710231718211A0032270936021606),
    .INIT_11(256'h09151F280B0B1E1F1C03261554080139341F093340420205041B170F12270423),
    .INIT_12(256'h1E0D081212072017050D000918202B3E3A1403170503052343100A1B22210910),
    .INIT_13(256'h3E070B2130140107160D0A1A150914060A34420004030604191D074D10060927),
    .INIT_14(256'h3D50471A302522071B32492A1B35181D0C0E090C0F0A180A05000A041F2D3230),
    .INIT_15(256'h2F00020716252B1201092F1B1D2A28142A210004070F0D4700183F210302030C),
    .INIT_16(256'h051A6D0406010803060D4C52390E18041221150C1E1D1E0F140F011345191A06),
    .INIT_17(256'h49032135291B0B0208040900080407010C3B03011E2F698A43164B1504220217),
    .INIT_18(256'h0000000000000000000000000000000B020805033836121D520F144148331513),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_785x450_sub_000000_351 (
    .addra({addra,3'b111}),
    .clka(clka),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa(doa[359:351]));
  // address_offset=0;data_offset=360;depth=785;width=9;num_section=1;width_per_section=9;section_size=450;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hB00206A9430000116901004451904780E5217C000020144019E21EE4684A6935),
    .INITP_01(256'h02022018000680804DFF0004F9C0CC9BF07EEFF11FFEF0E7FFB115FEFE217DE9),
    .INITP_02(256'h002D2181D5585D0C21092AC328CEA84388C48108206A123202AE630010627074),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000007500),
    .INIT_00(256'h00030202010100050703030002020102060C0C040C040605030301060608022D),
    .INIT_01(256'h10020D0701030003030603091200040F0B091E05421A0D090F08050509010203),
    .INIT_02(256'h15061125330C101425010700030820541119001D1F02073427275A455D524305),
    .INIT_03(256'h1A090A2B0F0C00133B2306483B0806023D0B066712033764453B2B31000B4941),
    .INIT_04(256'h04100324001909280108320A003E2D1D2F0E0133270B06170A04100511130709),
    .INIT_05(256'h0A04051617040D1614192C1520091F0415634C5F16100427101F0025060D040C),
    .INIT_06(256'h6209061016052101061F090F1E213238161B171C130E326C1836060E020B1808),
    .INIT_07(256'h2C15051E482A0B112E19050012020314321A2D0E0C0C0E0519070816342A0006),
    .INIT_08(256'h0C13233D3B06081E551006040D030E11070F01180412012F17081B1B05001429),
    .INIT_09(256'h4B7B5D554345223554010A03063D181C27080A0400051205382C4E5832232C02),
    .INIT_0A(256'h002D3119157E71977E6B4135500703394C6B21370D150003171D13050B103670),
    .INIT_0B(256'h1706142303313E321A1B454F5F353F1015130C01162C19482004151900010313),
    .INIT_0C(256'h1B18151C070C000B1A202833303F1204092804470E02130710311B0A3102180A),
    .INIT_0D(256'h231C4D2E2B15111419100E0A22120E01273F08212D190C040D09112050142E2D),
    .INIT_0E(256'h21150D3B353844250310050A07051101030C1211020C1F0E0C49251723180037),
    .INIT_0F(256'h0C07236A120C28270F69110A040508041010070B0005070B09101D01150F2927),
    .INIT_10(256'h16030103211816510C42065D5C3401121E071E0F011A0408061219040A070F15),
    .INIT_11(256'h2B2A080C07240F0502050A56034A032A3713112D11190F0701120A1B20260713),
    .INIT_12(256'h011007001426101023220A1F0A003A067913000A1D010706081A0205110F0333),
    .INIT_13(256'h33181628031B19051D040713031900070B0E240B76030202152F220708090B00),
    .INIT_14(256'h2A140E11111B0C0E3B162A2007060E1D040A1A2305012B0F3405090409271805),
    .INIT_15(256'h0C020B01100F3003043010020F051118131C1111070C05210C22096527010102),
    .INIT_16(256'h15072804010702030D090908181D221E3817250B0B04000C0D3512031D130841),
    .INIT_17(256'h60440C132A0005000105010006030A0E311D122D38573E1A300B1E28381F2A4D),
    .INIT_18(256'h0000000000000000000000000000000006060401070C00020008010700080A68),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_785x450_sub_000000_360 (
    .addra({addra,3'b111}),
    .clka(clka),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa(doa[368:360]));
  // address_offset=0;data_offset=369;depth=785;width=9;num_section=1;width_per_section=9;section_size=450;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h08001FCB63F9FCB7FFEBC9FFFBBC13F3EFD0F3ECCC77FFDF482B0C1301AC8D0A),
    .INITP_01(256'hF51D5E2337EFE1957F788865BD02211BD02A417F00E000F0665000327800036C),
    .INITP_02(256'h00434BDFCA173FFEE42040E200E1A8A0869BA01873BB00CFFC323E9B3513C383),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000012190),
    .INIT_00(256'h0A0102060005020206000400030101060100090A070502050006040302000646),
    .INIT_01(256'h00084D570E0003030300020011000509041F262F171311140502001107020204),
    .INIT_02(256'h570F0134040548550901010101020B124043453A2A1513573D081144473B0703),
    .INIT_03(256'h131913068660734E38203C0D0E00000004043C0D6D1D0275332A033D28074D25),
    .INIT_04(256'h6A3E041C012D0E14380F27605507445C0B00024E081B224D4817203F1C341033),
    .INIT_05(256'h30123B39361B395E280C1B0B0414041D2E485D630601074611324665592A336C),
    .INIT_06(256'h31291F313F39164613081B281A09010718302F1E6448652D174D012902292D1C),
    .INIT_07(256'h2C6E043F021B3A3506311819243B33200803021C1A37342B6F1D3D0F145B5714),
    .INIT_08(256'h0B563218365108304422410E2B120750696151442B052F1903121E1A34401819),
    .INIT_09(256'h080C0315093D31213456000C43566220283A35494B2D2E35341A15041C040511),
    .INIT_0A(256'h1B1718110D3407130C155C1B1000046F3B1A6D62471324170F14110B0810000D),
    .INIT_0B(256'h3509042410261B0A11160205101A4010350516666B2F0F200D2A120A491E3A1B),
    .INIT_0C(256'h1C18102D15030907021205050A0D0D04022A0630450003082B3B493D2110260B),
    .INIT_0D(256'h201C37273E08110D0A16291A12052D0905111706011B1D14291104033A2D2733),
    .INIT_0E(256'h1D0002194F014A542726240903260B1B1C17021B1E13040F1E21000E270E0527),
    .INIT_0F(256'h052C072E4D024E115C6E1704172A0D06151202020629031427060A0423211915),
    .INIT_10(256'h0805130118201405575509156F122C132D3B020004000E280F090B020C110510),
    .INIT_11(256'h201F10180A081327350427433D0506281E08150B464304011D020013280E0526),
    .INIT_12(256'h0C193A0B04110208100F040A0B08505D371110153D5D641E172D130A08140E18),
    .INIT_13(256'h1C130609151D0705060E010505160D2005172F1F48080D000A543A1837142C1E),
    .INIT_14(256'h34134D1606071F0A0C0D011403070A10071F050B182B37321D070405242A0C44),
    .INIT_15(256'h04040600181447142F240114031000100A150D001F061D015E08331801060505),
    .INIT_16(256'h49280010040202040105043E120A1E220B23041D0F2307041C30341F2E4E3233),
    .INIT_17(256'h6B1B1E172A291500030400000409463E0004210A1A000B075F0909343B101916),
    .INIT_18(256'h00000000000000000000000000000006040105190C3D17682C43231B323A015A),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_785x450_sub_000000_369 (
    .addra({addra,3'b111}),
    .clka(clka),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa(doa[377:369]));
  // address_offset=0;data_offset=378;depth=785;width=9;num_section=1;width_per_section=9;section_size=450;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h78F0FF8537FF41F07FF05407E7E409CC001C3300B0E0BE0D839F9DF63974EA56),
    .INITP_01(256'h56BFE000423C00860FC100C31E105C74FC28BFC3FA471A9E54109BDDC70B0DFE),
    .INITP_02(256'h03549F80D41C3BCD00001BD980017C40002F820006BC325001863F1044EB7F00),
    .INITP_03(256'h00000000000000000000000000000000000000000000000000000000000154F8),
    .INIT_00(256'h00050104050200060002020702070100040E060A01000302020C050401030423),
    .INIT_01(256'h0F020A3200020607020401221C22432A12133D3E120C04062812140103030906),
    .INIT_02(256'h083E3D50282849402D0201050704290A5003243D121B1A1946266A022009072E),
    .INIT_03(256'h081C3A3E4028089281600A31370202072924345F062A300E030E2E1E3D4C3515),
    .INIT_04(256'h2811140509241A17061D1C10061C4931000A020914434B09240304090B012525),
    .INIT_05(256'h12230227071A110B0C1C2706230503010D02295A0405000E425A0118170D1F24),
    .INIT_06(256'h0F3C112B011C1520060C0A07061C420B0B060A0F152D410B034C033734450513),
    .INIT_07(256'h2E6C02150E4F2F0A1E160E0B05071B1A07112A34281C29142902312F0842462A),
    .INIT_08(256'h03140326092F0B4103313D030C0A0A0106171E001F1D0E29181D160816281C30),
    .INIT_09(256'h070F060B00181F3918600563120C2F1A142001020517070F2028130C201F0003),
    .INIT_0A(256'h416E460506230C030B041F440804026A39520313130C0E1A0E220A0D3855081F),
    .INIT_0B(256'h090D2430222806161B0E0C08020A0A08480F055D152843401012150B000C0C3F),
    .INIT_0C(256'h1331221A08151204101B07020D20190E1E0622074301080B073C371718032920),
    .INIT_0D(256'h6A314D020701091B2F1D01132B1D240C25362421082A2B650E0C071795361102),
    .INIT_0E(256'h3A0B003C522C19062E0C0C050A14080624223A1736080F09070F34490A03072D),
    .INIT_0F(256'h40013001181004542E004225040F60281C1C0300002633272C031C040209251D),
    .INIT_10(256'h290D00100204130B34170B4F3D5C170A01163D0E293E0504090F394530131916),
    .INIT_11(256'h0215102319190722091B264C4A1E0427194D1C060D1E1E0D040510050C322638),
    .INIT_12(256'h132E171D060D1A0A101017090B07462B5A0C1422030418140603012508202105),
    .INIT_13(256'h1900161E1213242119150A0F0F051A261A01131C64000B066849302714132630),
    .INIT_14(256'h1C2D11245158280D3220233D331212040B302D6B300F08200B0200031A415D41),
    .INIT_15(256'h2C060702071F3A080F15491934242A131E0002050303326D582F203201070602),
    .INIT_16(256'h0C381402060C01000A09111331081E0F1A0B051212002418270A190D06420C27),
    .INIT_17(256'h513F28311C01050202070B03030A153B2F15101F321C2621221A1E041407513F),
    .INIT_18(256'h0000000000000000000000000000000A00010616121911372E463F3F191E4643),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_785x450_sub_000000_378 (
    .addra({addra,3'b111}),
    .clka(clka),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa(doa[386:378]));
  // address_offset=0;data_offset=387;depth=785;width=9;num_section=1;width_per_section=9;section_size=450;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hB081EE1F1000E370C27FF77B3D1AF1BF991CF2EFFD37819FB65FF67F300A67C8),
    .INITP_01(256'h05590E005181801E7C8E106DC132DEDE0D6FFBE3FDF5FFFDF34FFFFEFE530EF1),
    .INITP_02(256'h45AC10000520301E00091FFE08F4FDC897FFDD801BF118007F06C006804E8060),
    .INITP_03(256'h000000000000000000000000000000000000000000000000000000000000C8EC),
    .INIT_00(256'h05000408070A02000900030A0200060303100B11070106090309050507010800),
    .INIT_01(256'h0202483104010807030604231A224036183431551230011B041B140A0E090105),
    .INIT_02(256'h4D3C42110B3C1A440206040600034B1C0D022E431E451A3B0E3909373B46462D),
    .INIT_03(256'h0A040C0A05081D0A181512072301010001541D24281B14070A412A0120110942),
    .INIT_04(256'h240B042120050712041D0916164A2124260403011F28004A265106210B25321B),
    .INIT_05(256'h0B130E1F2A160310030F0204120E110F1118182C2A07050D0F3A3E3308190B07),
    .INIT_06(256'h5229000406162716070C17160F082D1A0915130B2B2217280C100F276544031A),
    .INIT_07(256'h46090F08004624100126191F1B321101070507121B2208081624096E380B6301),
    .INIT_08(256'h060A13390A040824111C0217112B08101D1701032F110F09070A080D01251657),
    .INIT_09(256'h1401050819022C463B59032233101F35320530220A253C2C512A03150E0C0700),
    .INIT_0A(256'h15130F2C0F17011E15100627490503022C2D3E2226313D151635222117220E1F),
    .INIT_0B(256'h064F41050B0107160B071B022E27201F0F07030A29120A1C0E2809070B140411),
    .INIT_0C(256'h060C2110082A44090D0C0E1719011405121619032D03040665210D221B0B0700),
    .INIT_0D(256'h690A11150E06060F040E08031C020C1C23070106080F2A4407110F01210F1515),
    .INIT_0E(256'h231704451B0D213015200A0F1D2D12041F000311301E0E0F2C160C021A140704),
    .INIT_0F(256'h35240B250B0B094F120B182A072B17012B3823191216071C3721272D3519040C),
    .INIT_10(256'h13001F17233724331651081C294E05010C2921161B352214100D0300001C102E),
    .INIT_11(256'h021D2F40332216031C3F290E1C56030E53260E280F2C00222910221F0A201C05),
    .INIT_12(256'h1D190B1D1300173624211D0D104D250E1D04020243433E1F09161D072C241D07),
    .INIT_13(256'h121C2B040A090622070B1D1B142430222B171622140507026F575B18102C2D13),
    .INIT_14(256'h0F49873E081D0F08130D17170A1B0C0A01314A0E07180B0A4302040155708508),
    .INIT_15(256'h19010800040F39562E28111804110812020E06031B171A12285587361C010908),
    .INIT_16(256'h5578580802040307051523144041330E3A10011C1A3A311C08110A1E081C2E0E),
    .INIT_17(256'h040E272312040501050B0B0105032636646019320D2F23304B2752407199650E),
    .INIT_18(256'h000000000000000000000000000000060A0302131200013407552405070A0813),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_785x450_sub_000000_387 (
    .addra({addra,3'b111}),
    .clka(clka),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa(doa[395:387]));
  // address_offset=0;data_offset=396;depth=785;width=9;num_section=1;width_per_section=9;section_size=450;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h00478C02DC39842C8998923DE08F803C55ECC306539933F9FB077F3F2C370148),
    .INITP_01(256'h137B0B801F70004924004FBBA007A221024220B024A10F80004C010F0C2010D0),
    .INITP_02(256'hC3B0300036FE00014FC5EE009C7EFD7B3A83D3FFF005FC9F74EFFCC7D8F788BE),
    .INITP_03(256'h000000000000000000000000000000000000000000000000000000000001A000),
    .INIT_00(256'h001009040507060202020504040101010105020600080D03010804040702030D),
    .INIT_01(256'h0A0E3B430202030801070402020B17110B22406A0732130D2101050D0E060203),
    .INIT_02(256'h04284A142E56634D2A000202040117170F0B2B3F2E3811312C590A0D33111731),
    .INIT_03(256'h18030B05081E0A071E020F312F0500042A0F185208110D030C01001A02353003),
    .INIT_04(256'h1D0C01012B233700210507300D0710341305031431371C05241B020F04091710),
    .INIT_05(256'h1E05170D180600011223190C0D2A101E0E0431031D080220081A05222C05000C),
    .INIT_06(256'h120C0A0B14100A0609091E0E18191C011D021A101701392B485E061E1D090F2D),
    .INIT_07(256'h3B470D243115290003080B1E1C07101A20221B2D170D2320191A343E3A335F1B),
    .INIT_08(256'h0A0A2466261315150C31032C12322A0E02250306040C33212C170215161A133D),
    .INIT_09(256'h222922120937007C3E5C05151212203517012207130D110A181E220A04071017),
    .INIT_0A(256'h1A0A080E180C222407471F434A070207373E11000119151E020B17121C0C2A1F),
    .INIT_0B(256'h0218352F22210F0C040A1307041F261E1C191731051506020F0516190213292D),
    .INIT_0C(256'h0F0C010C142F25190B1C061711100C051A04391204200F10002B070300040A0A),
    .INIT_0D(256'h100538072210121120303135220C0017101708000F200A041B150E096F1A2E17),
    .INIT_0E(256'h04100B4E201515050B0B0F01322B272623170B0D14200B1917060A1215080C1B),
    .INIT_0F(256'h1D12070741120A5536101C18160E1511081F2005011111081A0E0E220D0C1803),
    .INIT_10(256'h0E0F09191121111A201E0D27246735210A102006150616160C140A0418280513),
    .INIT_11(256'h16061C0F0418060021060118384E033A45880A2D0E0106130F06040A09130D27),
    .INIT_12(256'h1C011F130E0F0518151A220C0A0C0B12100C0E0F35290306080D001527422909),
    .INIT_13(256'h251901031314070E0207161D210611091B2503102B0411016C594919010B1D0B),
    .INIT_14(256'h57080306120911292A040505130D270609040B0C4317130D3A0408047E04362C),
    .INIT_15(256'h1202010220486B051937342200311F09220F2706111805070B01333440050000),
    .INIT_16(256'h3A2A3F020B050500080C5C524C26024955476C4206080E2A6502121108631A05),
    .INIT_17(256'h05010000011004040309080600051A10404A1A19516B2E09574D512331165C4A),
    .INIT_18(256'h0000000000000000000000000000000302060412353D1D062F691B1D58331220),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_785x450_sub_000000_396 (
    .addra({addra,3'b111}),
    .clka(clka),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa(doa[404:396]));
  // address_offset=0;data_offset=405;depth=785;width=9;num_section=1;width_per_section=9;section_size=450;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hF68E65FF1E8146E1B0765BA00E6A33C000261C810012CC079F27FFFF2A0E8517),
    .INITP_01(256'h429CFFF60417FFD079FFFD345E7E6B4217C0C414424C72066D5F08753BD7CE01),
    .INITP_02(256'hFE67DFFF0C6C139F20B37AE94B0017260031F945600B4C51012C6D7000897F70),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000012FFF),
    .INIT_00(256'h070004080500030000070702080701010C0501010501000D0A0600020209090E),
    .INIT_01(256'h0C07020F030303010001020202090F130A3D120A1E2F4A4A3513080F03020602),
    .INIT_02(256'h2A0723251507343C2F03030200010725171B043236200E2023693D610A3D2606),
    .INIT_03(256'h181005040928263B591D2B5D3A010508363B2E25153C340B0213262F3E1D031C),
    .INIT_04(256'h28020507070C080C0A2D120C15133058260309031F00031F122F090E1021171F),
    .INIT_05(256'h020622081104050F06132C1011060F0723020021050201052604373222030917),
    .INIT_06(256'h1F140B0F21030F190D0C1C0F29110A020F0F1A050D1A1F12073A010219320A23),
    .INIT_07(256'h803F070E3611101308070906090C03170E170905120C1B0F1B36503E5B603F0E),
    .INIT_08(256'h0A29082B720A0325201C2F010B1711030409241D192E09001616231E1019045D),
    .INIT_09(256'h1E2919020A092B17030801010F300A0F0515010301080D160621120701182106),
    .INIT_0A(256'h0F0B05001E0905190E071E1F191802431656120E0D1E04051F0F070D1B091E00),
    .INIT_0B(256'h0107000718240902050B18321C1D04194F1316116F59052105150B090C0F160D),
    .INIT_0C(256'h230208030B1302060D3004041D190608002F02080F0705096214140E0D1B0901),
    .INIT_0D(256'h77151B15111404161826090A0F1B190D0224594E1F5813435C0A030E7D251221),
    .INIT_0E(256'h42190014971823001C23050601241C03111E46454D7268583540030A6D17061B),
    .INIT_0F(256'h29100559341806290C2F1A1805010707100B3A202D314D56693D220E0C2D1032),
    .INIT_10(256'h243E2B141C2B00812B05121E11050A0E0B011704050D101803111D0D00240B1E),
    .INIT_11(256'h182F4B3B353623031A211C632206001404190A1611070C1712150C1102475639),
    .INIT_12(256'h0F060907141E231B331D232319041C1D0C0E1620073F111D200A061B00100607),
    .INIT_13(256'h030A051B170C0607261010041605191E1B0F372D07121C032829251D130A1412),
    .INIT_14(256'h451F33220919040329262303070D02211D1E09190522521B400109034A201563),
    .INIT_15(256'h040203051131463113151E11214301071D0305130207061132331C2211030004),
    .INIT_16(256'h002B3A180401040002010B282728300D0A2B1B2E0A1B0A334A000A172710092A),
    .INIT_17(256'h2E50442F20321B00030405050306012A5B2401833A331E69282538332D435253),
    .INIT_18(256'h0000000000000000000000000000000404000403070D1B3D6168523D4339285E),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_785x450_sub_000000_405 (
    .addra({addra,3'b111}),
    .clka(clka),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa(doa[413:405]));
  // address_offset=0;data_offset=414;depth=785;width=9;num_section=1;width_per_section=9;section_size=450;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h19B41B95DDE739179C7FB1EE07F1FF32DF1DFDD24F6F69A20E200000166A0B39),
    .INITP_01(256'hB1F030031007F83941EFE5380DF893C7FFC10C17F110F93E0B0B3B80C0B87021),
    .INITP_02(256'h384139F013FB9038AE189E12A904E7B9881FF85491FFC9E0788BDC040ABF8180),
    .INITP_03(256'h000000000000000000000000000000000000000000000000000000000001A000),
    .INIT_00(256'h05040205000409070807020509030203010C0808030005040102010206000305),
    .INIT_01(256'h1908320E010103000307091316172E220A36151B151F3B021A1A121104010506),
    .INIT_02(256'h2235054A42093C01160207030906223C0F0E021C4B0927090A01162731010341),
    .INIT_03(256'h0C060B091A191F2C080983050201070232335B1D294116083112032337261817),
    .INIT_04(256'h1714031201132007170501210517110A100405045A55781B1912090D0A0E0611),
    .INIT_05(256'h32001220212201130D06041B012812241C01080A030202022033310227200E1C),
    .INIT_06(256'h6C2E100416080516050A1F110A0C150C0105180D0400060D2E0E002D063B241C),
    .INIT_07(256'h8019033B3314103215191718071B0809140D1E18140006300622180B99015A5B),
    .INIT_08(256'h011315465B2901266F0D051B18120E0B090D1A260C260E0D01000E061B212F07),
    .INIT_09(256'h2516180C1C090D0B8B45012E50302C210F050704050B071E12331D1B15310B14),
    .INIT_0A(256'h102D1415020F1C17263A1F567B220B264C2A070D0D09070418070A0E2601040F),
    .INIT_0B(256'h241F0B20121E32360702190F251039644228000241321E3C03110B0B00071415),
    .INIT_0C(256'h3F10190A280D051D2914022B2601090B05150B844727163584062C3E0002160D),
    .INIT_0D(256'h0E0C2E4E483A280304122204353C12301F1A06150710033D362206181D024142),
    .INIT_0E(256'h0612084D1F153D1538123C0E2415400A1A180C0609052F25353D0322141A1635),
    .INIT_0F(256'h0201152D35040963191D1B0C1D0A0E2E1D2A150F1C090E122D213E5236291626),
    .INIT_10(256'h1F222F12071A2522071A03668E163A2606170B2820401704070E23304140381B),
    .INIT_11(256'h2A0601051C2501001706000C3931032E59281023150D051B16302911072B2625),
    .INIT_12(256'h05182B082F050B11241C0428250E213B5D260000462C510D0224041504242514),
    .INIT_13(256'h0208080B03021811040E261E1A02132F0E205E4944070A02380C451210081606),
    .INIT_14(256'h4C0E1408221D080B010C06160612020F1B2A1E053F0A57401D0401010C2B0803),
    .INIT_15(256'h05000404160C1A4F282B1B150844312318001F0817181D1F4A5E331F23010100),
    .INIT_16(256'h1E283E02060607070708383C0A0A2D1D13032722351E222738300B4A39091E06),
    .INIT_17(256'h64251C25090F000703010B030005010E6C3A121A040E102E2E3A2D2A1956311F),
    .INIT_18(256'h000000000000000000000000000000040201080F5A8774567E8C343A84542A6C),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_785x450_sub_000000_414 (
    .addra({addra,3'b111}),
    .clka(clka),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa(doa[422:414]));
  // address_offset=0;data_offset=423;depth=785;width=9;num_section=1;width_per_section=9;section_size=450;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hCCC000FB9801061FCCF000DDC0083C41E7319C788050FA4127E71AE2401D0135),
    .INITP_01(256'h0EBEA0037C01903C80003FE4321FF4D3F3FF2F3DFFBAFFFE0187F1E00CEE2050),
    .INITP_02(256'h0018F630F23B8D04A15AF9D59FCBA5A8181DA300417A33A77D2770A044622910),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000016D80),
    .INIT_00(256'h010408070405010206000D01040C0A01020A000809050A070A0003020302020A),
    .INIT_01(256'h06040501060106030707050100060A09080F104D34002A090F1101010A060609),
    .INIT_02(256'h0446270779350219120500040008203427236162010C0425150F0B0335344802),
    .INIT_03(256'h14060C0F01293B071B001C060F00010208020A382C1A00510A411C1017001622),
    .INIT_04(256'h141A1C070611050E1E333409051A3306130103010437250404151E151E04021C),
    .INIT_05(256'h0302261C170D1F010C190B074229030A0024233D000C02031B2D051D3403020E),
    .INIT_06(256'h261429070E062111011A0E00010B0A071313030300241C7B182401115F270524),
    .INIT_07(256'h052503062803002E061C0F0B160D020C2F2930280C0D0D0B330C071B2D1F050E),
    .INIT_08(256'h203421110E2D022F2B54222E033A020E0A13090600023F120809020709380807),
    .INIT_09(256'h0403401B244329044602002900271D4D1A16190A041B06092A342D041B1D201C),
    .INIT_0A(256'h2B868F9B734D1A1A1D27053456040303534C5E2F110A110E1C05150D29685103),
    .INIT_0B(256'h141A070214231E657A8F8366583B7B50200D19040E3C241201021D12140A0214),
    .INIT_0C(256'h0111110405220907132E29010F4289A2ACFFA6541511051D1310141407121710),
    .INIT_0D(256'h060F42522A240C02061609150E1B0C1F21031930619E644A07130A1842261202),
    .INIT_0E(256'h07120508201A033E0C180C310D0C050B0632150102130D1735023F3D1012080E),
    .INIT_0F(256'h05342857261002460A1F170A191D0C14180F0B00171C260A23151920292A1104),
    .INIT_10(256'h030A0805030433420A1113375F1E29110700091F0B0E0F0B0916290A000D1126),
    .INIT_11(256'h070A220D0C030D06091E123A4F070806481623080C080A281C060A0512080B22),
    .INIT_12(256'h18010C06140D070E0B0A0F0F09262D012F190B123B2C0A110F1C0B0C0E0F0C06),
    .INIT_13(256'h07260707070A1D0C070B0804150217011109120F440006041550322C0F2A1124),
    .INIT_14(256'h06430C072725162E1D3F001E021C06011B160E192A0100092A070F050D380515),
    .INIT_15(256'h2600010C090750200F0A0E081008171C060A0C13132404070E06892F23050706),
    .INIT_16(256'h1F3F2802000203000D012E450103032E0D0A2A2B0B2D1C2228422B32021E0473),
    .INIT_17(256'h695A210B130400040407000505100B024B642408033823715D080D19130C185F),
    .INIT_18(256'h000000000000000000000000000000050A0207044336012D250A5D7156364B7B),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_785x450_sub_000000_423 (
    .addra({addra,3'b111}),
    .clka(clka),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa(doa[431:423]));
  // address_offset=0;data_offset=432;depth=785;width=9;num_section=1;width_per_section=9;section_size=450;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h00508461840A765C000A053FC3F1B12C7EE90913F8FCF7FF821F95FC4C2E90D8),
    .INITP_01(256'h160F8F21FED8D41D812E01BB22801BA32900B42AEC0103B002083F0A0401B0F6),
    .INITP_02(256'h0650310A00FFCE7C6EDD3D8487F059A17F005677E800FFFE058BD22570B55866),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000015840),
    .INIT_00(256'h0504020101020604000A020101020300030800020200000009080A0104050616),
    .INIT_01(256'h11032340050404060B00041319153A320929212C0B03000F2415170D10050B03),
    .INIT_02(256'h072B3C822B1B433C340A0308080A11211949352E2B1B6B76606A18748E815F24),
    .INIT_03(256'h040A073322162A0F66252E02300305020D290B3B0227092303190A1F3E001F07),
    .INIT_04(256'h02030000160E05051F0C11071F271A2E3C07071333631F1719200D0E06160A22),
    .INIT_05(256'h1B0F1D260D231016000F10090A0001000F3314003C05000B193D1C420B0D0309),
    .INIT_06(256'h2727453B0A16081E2733110B290B011B001C1A15180E41283A08022B192D031B),
    .INIT_07(256'h493D032C0F2F640F130C1A0A1E101F1B111213270E0A0209262A2041980A5C27),
    .INIT_08(256'h1E30121C251F041100585223072C330A2711100B021115110C2A1C070811440B),
    .INIT_09(256'h0900303528190B77535807070500321B4A09081D060C0A0D1507130D0705200E),
    .INIT_0A(256'h0307040B0602143D2848356B3200054050352C15220622310A0C070113162409),
    .INIT_0B(256'h120502080C0A060C12022A2E1E215950450F203C09180D1B0B0B110502070902),
    .INIT_0C(256'h0E29120026121807111304121504162917480541421305161B0E2C02331B090C),
    .INIT_0D(256'h350C1520220D02080F1A060A12040406100C141C142432583B0A140B5D171D03),
    .INIT_0E(256'h090B010B442235000E0928120A30100401170810010D130A1A072E4249020E18),
    .INIT_0F(256'h1A1D211621180A41320B0400211201230137230F180F130605061C140B243922),
    .INIT_10(256'h0C02040B0524161D0D0E102B084E090205160305011B2816020D05100220090A),
    .INIT_11(256'h081603171C010B14180C07032D48063C1C760617080B0107131C07040F1D0909),
    .INIT_12(256'h350425050811000C0D1714060D1D19026F0E1313112B2C2D140809091E1A1D00),
    .INIT_13(256'h2F182D1D3F1814030913221C1D060A061C0C070214080D03592C420B0D144827),
    .INIT_14(256'h4B44061B0E0717152C1D1D0E091004121814120A1100051C2804010914200128),
    .INIT_15(256'h1D0108002D3B38100248263A185305030424031C2504050109154301220C0205),
    .INIT_16(256'h0C1E601906050C05090D43271E190D1F2D053626090F1C2523381D043C3B063F),
    .INIT_17(256'h271417231F0B0A000602040705021737631E0924282602195022651017170908),
    .INIT_18(256'h000000000000000000000000000000020004011C02061A551C3410231B08323D),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_785x450_sub_000000_432 (
    .addra({addra,3'b111}),
    .clka(clka),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa(doa[440:432]));
  // address_offset=0;data_offset=441;depth=785;width=9;num_section=1;width_per_section=9;section_size=450;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hDFEEE539D99993B770BA9CEFFBBFC0FCB7FC15D800C8C840CCA411C722226590),
    .INITP_01(256'h8CFFC039E268629C8E0861C4F0825D53006363A00BF6B880CF31FC21345DE45A),
    .INITP_02(256'h06650006EA039E40306AFEC957FFC7B5BFFFF83FFFE8B1FFFFCF69E4F8ACEC03),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000003040),
    .INIT_00(256'h070A030A0506020403000505000B0202000F0D000707010306050B0902030700),
    .INIT_01(256'h01023E440203000109000913080705120336401F083E030E2D0D021516020108),
    .INIT_02(256'h6E53730520424E4C2103040802090F06484803180D224B43193F1D553B1C332F),
    .INIT_03(256'h19082337290635594117621D2707020B210F4B2C3C1B1C655A040D050303107B),
    .INIT_04(256'h355E4B111C062F4C200530302B2E0C4F2D01014D0E1C23082141300C0E073A03),
    .INIT_05(256'h0F02301B11100C000327141621161805160C1474370D094F1856041B05571A0E),
    .INIT_06(256'h04181C0F3C030A1F03180028040002011722274517101D5C562E031B0D3F0F19),
    .INIT_07(256'h372205121F2D02100C1B0804170715000D1B0D1D13011E221814AA803F611D25),
    .INIT_08(256'h1210221E2746011B16510030052001071B0D1404170C15141E07250C0721663D),
    .INIT_09(256'h0B15191A1D211B460853012803340B0E130A09082B0F270715120A041B130004),
    .INIT_0A(256'h3A0B080D0A00050E0D1620474B0609436621141C220318090412242510161710),
    .INIT_0B(256'h2825282038541F07171E01160D0C25364A0C135C09333E3403020A132D1F3D2E),
    .INIT_0C(256'h041B1D054C0F1E0A0227231E2418140E2D11070D1018000E180630200B083B04),
    .INIT_0D(256'h070F2D03011B38293A441D171E031C1215042C071D28042A0D06000941031604),
    .INIT_0E(256'h0F0A0867101F030824041412052A422408060B121D0403260A173226231D052C),
    .INIT_0F(256'h281657101A1B52902A060E140C0D050709072E37071D2827221608281A3D3417),
    .INIT_10(256'h051125203708404B0A2A0752250B0B1410060B15081A0A2D2B1A1C331003032B),
    .INIT_11(256'h170E0E0F2D043D13212D105D5823050710211D201D0A0003020B180C2D070E15),
    .INIT_12(256'h0C6343604437273C293036041C0213335F060812004F1C27232D2D302C1D4339),
    .INIT_13(256'h0820083729584C2A23452C2E1720090905360F084804000961301E663E273624),
    .INIT_14(256'h23240C2C001A0D4A3832202A1B1E1C2C071C0E30190D1F150E040A010A240912),
    .INIT_15(256'h1A0509061C0A891E0A051C02121919021424513D2629040B220D2F0810010308),
    .INIT_16(256'h031A011B09010300030C3A14284E012116172216040715280505114D5C373011),
    .INIT_17(256'h281A16090620100A0F040B0300070E02273C91541A001A44581507080008163A),
    .INIT_18(256'h000000000000000000000000000000060002010C0F1A1C4A521044456C18361C),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_785x450_sub_000000_441 (
    .addra({addra,3'b111}),
    .clka(clka),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa(doa[449:441]));

endmodule 

