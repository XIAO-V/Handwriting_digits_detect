// Verilog netlist created by TD v4.6.18154
// Fri Nov 13 14:37:04 2020

`timescale 1ns / 1ps
module rom_digit  // al_ip/word/result.v(14)
  (
  addra,
  clka,
  rsta,
  doa
  );

  input [12:0] addra;  // al_ip/word/result.v(18)
  input clka;  // al_ip/word/result.v(19)
  input rsta;  // al_ip/word/result.v(20)
  output [10:0] doa;  // al_ip/word/result.v(16)

  wire [0:1] addra_piped;
  wire  \inst_doa_mux_b0/B0_0 ;
  wire  \inst_doa_mux_b0/B0_1 ;
  wire  \inst_doa_mux_b1/B0_0 ;
  wire  \inst_doa_mux_b1/B0_1 ;
  wire  \inst_doa_mux_b10/B0_0 ;
  wire  \inst_doa_mux_b10/B0_1 ;
  wire  \inst_doa_mux_b2/B0_0 ;
  wire  \inst_doa_mux_b2/B0_1 ;
  wire  \inst_doa_mux_b3/B0_0 ;
  wire  \inst_doa_mux_b3/B0_1 ;
  wire  \inst_doa_mux_b4/B0_0 ;
  wire  \inst_doa_mux_b4/B0_1 ;
  wire  \inst_doa_mux_b5/B0_0 ;
  wire  \inst_doa_mux_b5/B0_1 ;
  wire  \inst_doa_mux_b6/B0_0 ;
  wire  \inst_doa_mux_b6/B0_1 ;
  wire  \inst_doa_mux_b7/B0_0 ;
  wire  \inst_doa_mux_b7/B0_1 ;
  wire  \inst_doa_mux_b8/B0_0 ;
  wire  \inst_doa_mux_b8/B0_1 ;
  wire  \inst_doa_mux_b9/B0_0 ;
  wire  \inst_doa_mux_b9/B0_1 ;
  wire \and_Naddra[11]_addra_o ;
  wire inst_doa_i0_000;
  wire inst_doa_i0_001;
  wire inst_doa_i0_002;
  wire inst_doa_i0_003;
  wire inst_doa_i0_004;
  wire inst_doa_i0_005;
  wire inst_doa_i0_006;
  wire inst_doa_i0_007;
  wire inst_doa_i0_008;
  wire inst_doa_i0_009;
  wire inst_doa_i0_010;
  wire inst_doa_i2_000;
  wire inst_doa_i2_001;
  wire inst_doa_i2_002;
  wire inst_doa_i2_003;
  wire inst_doa_i2_004;
  wire inst_doa_i2_005;
  wire inst_doa_i2_006;
  wire inst_doa_i2_007;
  wire inst_doa_i2_008;
  wire inst_doa_i2_009;
  wire inst_doa_i2_010;

  reg_sr_as_w1 addra_pipe_b0 (
    .clk(clka),
    .d(addra[11]),
    .en(1'b1),
    .reset(rsta),
    .set(1'b0),
    .q(addra_piped[0]));
  reg_sr_as_w1 addra_pipe_b1 (
    .clk(clka),
    .d(addra[12]),
    .en(1'b1),
    .reset(rsta),
    .set(1'b0),
    .q(addra_piped[1]));
  and \and_Naddra[11]_addra  (\and_Naddra[11]_addra_o , ~addra[11], addra[12]);
  EG_PHY_CONFIG #(
    .DONE_PERSISTN("ENABLE"),
    .INIT_PERSISTN("ENABLE"),
    .JTAG_PERSISTN("DISABLE"),
    .PROGRAMN_PERSISTN("DISABLE"))
    config_inst ();
  // address_offset=0;data_offset=0;depth=4096;width=8;num_section=1;width_per_section=8;section_size=11;working_depth=4096;working_width=8;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM32K #(
    .CLKBMUX("0"),
    .CSAMUX("INV"),
    .CSBMUX("0"),
    .DATA_WIDTH_A("8"),
    .DATA_WIDTH_B("8"),
    .INIT_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_04(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_05(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_06(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFEFAFAFAFAFAFBFBFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'hDFDFDFDFDFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0A(256'hFFFFFFDFDFDFDFDFDFDF9F9F9F9D989898DADADAD2D2D2D2D2D2D2DADADADBDB),
    .INIT_0B(256'h5252525253535B5F5F5F7F7F7F7F7F7F7F7F7FFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0C(256'hFFFF7F7F7F7F7F5F1F0F0F0F0F0F0F0E0A080800101012121212525252525252),
    .INIT_0D(256'h125252525252525252525353535F7F7F7F7F7F7F7F7F7FFFFFFFFFFFFFFFFFFF),
    .INIT_0E(256'hFFFFFFFFFFFF7F7F7F7F3F1F1F0F0F0F0F0E0A0A020000001010101012121212),
    .INIT_0F(256'h101212121212125252525252525252525353777F7F7F7F7F7F7F7FFFFFFFFFFF),
    .INIT_10(256'hFFFFFFFFFFFFFFFFFFFF7F7F7F3F3F1F1F0F0F0F0A0A02020200000000101010),
    .INIT_11(256'h001010101010101212121212125252525252525252537373777F7F7F7F7F7FFF),
    .INIT_12(256'h7F7F7FFFFFFFFFFFFFFFFFFFFFFF7F7F7F3F3F1F1F0F0F0A0A02020202000000),
    .INIT_13(256'h02000000000010101010101010121212121252525252525252527373737F7F7F),
    .INIT_14(256'h737B7F7F7F7F7FFFFFFFFFFFFFFFFFFFFFFF7F7F7F3F3F1F1F0F0A0A02020202),
    .INIT_15(256'h0202020202000000000010101010101010101012121212525252525252527273),
    .INIT_16(256'h52527272737B7B7F7F7F7FFFFFFFFFFFFFFFFFFFFFFF7F7F7F3F3F1F1F0A0A02),
    .INIT_17(256'h1A0A020202020202020000000000011515151515151515141416121252525252),
    .INIT_18(256'h1652525252527272737B7B7F7F7F7FFFFFFFFFFFFFFFFFFFFFFFFF7F7F3F3F1F),
    .INIT_19(256'h7F3F3F3B3A2222626262626262606060656565353D3D3D3D3D3D3D3D3D3C1C1E),
    .INIT_1A(256'hBDBD9C9C9C9EDED2D2D2D2F2F2FBFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7F),
    .INIT_1B(256'hFFFFFFFF7F3F3F3A7262626262E2E2E2E2E0E1E5E5EDEDEDFDFDBDBDBDBDBDBD),
    .INIT_1C(256'hBDBDBDBDBDBD9D9C9C9C9CDEDAD2D2F2F2FAFBFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1D(256'hFFFFFFFFFFFFFFFF7F3F7A7A7262626262E2E2E2E2E1E5E5EDEDEDEDFDFDFDFD),
    .INIT_1E(256'hEDFDFDFDFDBDBDBDBDBD9D9D9C9C9C9CDCDCDAF2F2FAFBFFFFFFFFFFFFFFFFFF),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFF7F7A72726262626262E2E2E2E5E5EDEDEDEDED),
    .INIT_20(256'hEDEDEDEDEDEDFDFDFDFDBDBDBDBD9D9D9D9C9C9C9CDCDCF8F0FAFAFFFFFFFFFF),
    .INIT_21(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFA7A72726262626262E2E2E7E5EDED),
    .INIT_22(256'hE7EDEDEDEDEDEDEDEDEDFDFFFFFDFDBDBDBD9D9D9D9D9C9C9CDCDCFCF8FAFAFF),
    .INIT_23(256'hFCFEFAFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFA7A7272626262626262E7),
    .INIT_24(256'h62626267E7EDEDEDEDEDEDEDEDEDEDFFFFFFFDFDBDBD9D9D9D9D9C9C9C9CDCFC),
    .INIT_25(256'h9C9CDCFCFCFEFEFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFAFA7272626262),
    .INIT_26(256'h7262626262626767EFEDEDFDEDEDEDEDEDEDEDFFFFFFFFFFFDBD9D9D9D9D9D9C),
    .INIT_27(256'h9D9D9D9C9C9C9CFCFCFEFEFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFAFA72),
    .INIT_28(256'hFAFAF2F272626262626267676FEDEDFDEDEDEDEDEDEDEDEFFFFFFFFFFFFF9D9D),
    .INIT_29(256'hFFFFDF9F9D9D9D9C9C9C9CBCFCFEFEFEFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_2A(256'hFFFFFFFFFAFAF2F272626262626367676FEDEDFDFDEDEDEDEDEDEDEFEFFFFFFF),
    .INIT_2B(256'hEFFFFFFFFFFFFF9F9F9F9D9D9C9C9CBCFCFEFEFEFEFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_2C(256'hFFFFFFFFFFFFFFFEFAFAF2F2F2626262626367676F6DEDFDFDEDEDEDEDEDEDEF),
    .INIT_2D(256'hEDEDEDEFEFEFFFFFFFFFFFDF9F9F9F9F9C9C9CBCFCFEFEFEFEFFFFFFFFFFFFFF),
    .INIT_2E(256'hFFFFFFFFFFFFFFFFFFFFFFFEFAFAF2F2F2626262626367676F6DEDFDFDFDEDED),
    .INIT_2F(256'hFDFDEDEDEDEDEDEFEFEFEFFFFFFFFFDF9F9F9F9F9E9E9EBCBCFEFEFEFEFEFFFF),
    .INIT_30(256'hFEFEFFFFFFFFFFFFFFFFFFFFFFFFFFFEFAFAF2F2F2E26262626367676F6D6DFD),
    .INIT_31(256'h6F6D6DFDFDFDFDEDEDEDEDEFEFEFEFFFFFFFFFDFDF9F9F9F9F9E9EBEBEFEFEFE),
    .INIT_32(256'hBEBEFEFEFEFEFFFFFFFFFFFFFFFFFFFFFFFFFFFEFAFAFAF2F2E2E26263636767),
    .INIT_33(256'h636367676F6D6D7DFDFDFDFDEDEDEDEFEFEFEFEFFFFFFFDFDF9F9F9F9F9E9EBE),
    .INIT_34(256'h9F9E9E9EBEBEFEFEFEFEFFFFFFFFFFFFFFFFFFFFFFFFFFFEFAFAFAF2F2E2E262),
    .INIT_35(256'hF2E2E2E2636367676F6D6D7DFDFDFDFDEDEDEDEFEFEFEFEFEFFFFFDFDF9F9F9F),
    .INIT_36(256'hDFDF9F9F9F9E9E9EBEBEFEFEFEFEFEFFFFFFFFFFFFFFFFFFFFFFFEFEFEFAFAF2),
    .INIT_37(256'hFEFAFAF2F2E2E2E2636367676F6D6D7D7DFDFDFDFDEDEDEFEFEFEFEFEFFFFFDF),
    .INIT_38(256'hEFEFFFDFDFDF9F9F9F9E9E9EBEBEBEFEFEFEFEFFFFFFFFFFFFFFFFFFFFFFFEFE),
    .INIT_39(256'hFFFFFEFEFEFAFAF2F2E2E2E2E3636767676D6D7D7D7DFDFDFDEDEDEFEFEFEFEF),
    .INIT_3A(256'hEFEFEFEFEFEFEFDFDFDF9F9F9F9F9E9EBEBEBEFEFEFEFEFFFFFFFFFFFFFFFFFF),
    .INIT_3B(256'hFFFFFFFFFFFFFEFEFEFAFAFAF2E2E2E3E3636367676D6D7D7D7DFDFDFDFDEDEF),
    .INIT_3C(256'hFDFDFDEFEFEFEFEFEFEFEFDFDFDFDF9F9F9F9E9EBEBEBEFEFEFEFEFFFFFFFFFF),
    .INIT_3D(256'hFFFFFFFFFFFFFFFFFFFFFEFEFEFAFAFAF2E2E2E3E3E36367676D6D7D7D7D7DFD),
    .INIT_3E(256'h7D7D7DFDFDFDFDEFEFEFEFEFEFEFEFCFDFDFDF9F9F9F9E9EBEBEBEFEFEFEFEFF),
    .INIT_3F(256'hFEFEFEFFFFFFFFFFFFFFFFFFFFFFFEFEFEFEFAFAFAE2E2E3E3E3636367656D7D),
    .INIT_40(256'h6765653D3D3D3D3DBDFDFDFFEFEFEFEFEFEFEFCFCFDFDF9F9F9F9E9EBEBEBEFE),
    .INIT_41(256'hBEBEBEBEFEFEFEFFFFFFFFFFFFFFFFFFFFFFFEFEFEFEFAFAFAE2E2E3E3E3E363),
    .INIT_42(256'hE3E3A323232525353D3D3D3DBD9D9D9F9FCFCFEFEFEFEFCFCFDFDF9F9F9F9E9E),
    .INIT_43(256'h9F9F9E9EBEBEBEBEFEFEFEFFFFFFFFFFFFFFFFFFFFFFFEFEFEFEFAFAFAEAE2E3),
    .INIT_44(256'hFAEAEAE3A3A3A3A323252515151D1D1D1D9D9D9F9F8F8F8FCFCFCFCFCFCFDF9F),
    .INIT_45(256'hCFCFCF9F9F9F9E9EBEBEBEBEFEFEFEFFFFFFFFFFFFFFFFFFFFFFFEFEFEFEFEFA),
    .INIT_46(256'hFEFEFEFAFAEAAAABA3A3A3A3030105151515151D1D9D9D9F9F9F8F8F8FCFCFCF),
    .INIT_47(256'h8F8F8FCFCFCFCFDF9F9F9E9EBEBEBEBEFEFEFEFFFFFFFFFFFFFFFFFFFFFEFEFE),
    .INIT_48(256'hFFFEFEFEFEFEFEFEBAAAAAABABA38383830101151515151515159D9F9F9F9F8F),
    .INIT_49(256'h9797978787878787C7C7C7C79F9F9E9EBEBEBEBEFEFEFEFEFFFFFFFFFFFFFFFF),
    .INIT_4A(256'hFFFFFFFFFFFEFEFEFEFEFEBEBEAAAAAB8B8B8B83830101111515151515159597),
    .INIT_4B(256'h151595979797979787878787C7C7C7C78F9F9E9EBEBEBEBEFEFEFEFEFFFFFFFF),
    .INIT_4C(256'hFFFFFFFFFFFFFFFFFFFEFEFEFEFEBEBEBEAAAA8B8B8B8B8B8B01011111151515),
    .INIT_4D(256'h1111151515151597979797979787878787C7C7C78F8F9E9EBEBEBEBEFEFEFEFE),
    .INIT_4E(256'hFEFEFEFEFFFFFFFFFFFFFFFFFFFEFEFEFEBEBEBEBE8E8A8B8B8B8B8B8B890911),
    .INIT_4F(256'h8B89095959515155555555D7D7D79797978787878787C7C78F8F9E9E9EBEBEBE),
    .INIT_50(256'hBEBEBEBEBEFEFEFEFFFFFFFFFFFFFFFFFFFEFEFEFEBEBEBE9E8E8E8B8B8B8B8B),
    .INIT_51(256'h8B8B8B8B8BC1C1515151515151557577F7F7F7F7B7B7A7A7A7A7A7E7AFAFAEBE),
    .INIT_52(256'hAFAFAEAEBEBEBEBEBEFEFEFEFFFFFFFFFFFFFFFFFFFEFEFEBEBEBEBE9E8E8E8F),
    .INIT_53(256'h9E8E8E8F8F8B83C3C3C1C1515151717171717577F7F7F7F7F7B7B7A7A7A7A7A7),
    .INIT_54(256'hA7A7A7A7AFAFAEAEAEBEBEBEBEFEFEFEFFFFFFFFFFFFFFFFFFFEFEBEBEBEBE9E),
    .INIT_55(256'hBEBE9E9E9E8E8E8F8787C3C3C3C1C1D1717171717171717777F7F7F7F7F7B7B7),
    .INIT_56(256'hF7F7F7B7A7A7A7A7AFAFAEAEAEBEBEBEBEFEFEFEFFFFFFFFFFFFFFFFFFFEFEBE),
    .INIT_57(256'hFFFEBEBEBEBE9E9E9E8E868787C7C7C3C3C1C1F1717171717171717373F7F7F7),
    .INIT_58(256'h7B7BFFFFFFFFFFFFBFAFAFAFAFAFAEAEAEAEBEBEBEFEFEFEFFFFFFFFFFFFFFFF),
    .INIT_59(256'hFFFFFFFFFFFEBEBEBE9E9E9E9E86868787C7C7C7C3E1E1F1717171717179797B),
    .INIT_5A(256'h7979797B7B7BFBFFFFFFFFFFFFBFAFAFAFAFAEAEAEAEAEBEBEFEFEFEFFFFFFFF),
    .INIT_5B(256'hFFFFFFFFFFFFFFFFFFFFBEBEBE9E9E9E96868687C7C7C7C7E7E5E1F1F1797979),
    .INIT_5C(256'hF97979797979797B7B7BFBFBFBFFFFFFFFFFAFAFAFAFAEAEAEAEAEAEBEFEFEFE),
    .INIT_5D(256'hAEFEFEFFFFFFFFFFFFFFFFFFFFBFBEBE9E9E9E96968686C7C7C7C7E7E7E5E5F9),
    .INIT_5E(256'hE7E5EDFDF9F979797979797B7B7B7BFBFBFBFFFFFFFFBFAFAFAFAEAEAEAEAEAE),
    .INIT_5F(256'hAEAEAEAEAEEEFEFFFFFFFFFFFFFFFFFFFFBFBEBE9E9E9696968686C7C7C7C7E7),
    .INIT_60(256'hC7C7E7E7E7EDEDFDFDFD79797979797B7B7B7BFBFBFBFBFFFFFFBFBFAFAFAEAE),
    .INIT_61(256'hBFAFAEAEAEAEAEAEAEEEFEFFFFFFFFFFFFFFFFFFFFBFBEBE9E9E9696968686C7),
    .INIT_62(256'h9686C6C7C7C7E7E7EFEDEDFDFDFD7D797979797B7B7B7B7BFBFBFBFBFBFFFFBF),
    .INIT_63(256'hFBFBFFBFBFBFAEAEAEAEAEAEEEEEEEFFFFFFFFFFFFFFFFFFFFBFBEBE9E969696),
    .INIT_64(256'h9E9696969686C6C7C7E7E7EFEFEDEDFDFDFDFD7D7D79797B7B7B7B7BFBFBFBFB),
    .INIT_65(256'hFBFBFBFBFBFBFBBFBFBFAEAEAEAEAEAEEEEEEEEFFFFFFFFFFFFFFFFFFFBFBEBE),
    .INIT_66(256'hBFBFBE9E969696969686C6C7C7E7EFEFEFEDEDFDFDFDFD7D7D7D797B7B7B7B7B),
    .INIT_67(256'h7B7B7B7B7BFBFBFBFBFBFBBBBFBFBEAEAEAEAEAEEEEEEEEFEFFFFFFFFFFFFFFF),
    .INIT_68(256'hFFFFFFFFBFBFBE9E969696969686C6C7C7E7EFEFEFEDEDFDFDFDFDFD7D7D7D7F),
    .INIT_69(256'h6D6D6D6F6F6B6B6B6BEBEBEBEBEBEBABABAEAEAEAEAEAEAEEEEEEEEFEFEFFFFF),
    .INIT_6A(256'hEFEFFFFFFFFFEFEFAFAFAE8E868686868686C6C6C7EFEFEFEFEDEDEDEDEDEDED),
    .INIT_6B(256'hEDEDEDED6D6D6D6F6F6F6B6B6B6BEBEBEBEBEBABABAAAEAEAEAEAEAEEEEEEEEF),
    .INIT_6C(256'hEEEEEEEFEFEFFFFFFFFFEFEFAFAFAF8E868686868686C6C6C7EFEFEFEFEDEDED),
    .INIT_6D(256'hEFEDEDEDEDEDEDEDED6D6D6F6F6F6F6F6B6BEBEBEBEBEBABABAAAAAEAEAEAEAE),
    .INIT_6E(256'hAEAEAEAEEEEEEFEFEFEFFFFFFFFFEFEFAFAFAF86868686868686C6C6C7EFEFEF),
    .INIT_6F(256'hC7EFEFEFEFEDEDEDEDEDEDEDED6D6D6F6F6F6F6F6F6BEBEBEBEBEBABABAAAAAA),
    .INIT_70(256'hABAAAAAAAAAEAEAEEEEEEFEFEFEFFFFFFFFFEFEFAFAFAF86868686868686C6C6),
    .INIT_71(256'h8686C6C6C7EFEFEFEFEDEDEDEDEDEDEDED6D6D6F6F6F6F6F6F6F6BEBEBEBEBAB),
    .INIT_72(256'hEBEBEBABAAAAAAAAAAAEAEEEEEEEEFEFEFEFFFFFFFFFEFEFAFAFAF8686868686),
    .INIT_73(256'h868686868686C6C6C6EFEFEFEFEDEDEDEDEDEDEDEDED6D6F6F6F6F6F6F6F6FEB),
    .INIT_74(256'h6F6F6FEFEBEBEBABAAAAAAAAAAAAAEEEEEEEEFEFEFEFFFFFFFFFEFEFEFAFAFA7),
    .INIT_75(256'hEFAFAFA7868686868686C6C6C6EFEFEFEFEDEDEDEDEDEDEDEDED6D6F6F6F6F6F),
    .INIT_76(256'h6F6F6F6F6F6F6F6FEFEBABABAAAAAAAAAAAAAAEEEEEFEFEFEFEFFFFFFFFFEFEF),
    .INIT_77(256'hFFFFEFEFEFAFAFAF868686868686C6C6C6CFEFEFEFEDEDEDEDEDEDEDEDED6D6F),
    .INIT_78(256'hFDFDFD7F7F7F7F7F7F7F7F7FFFFFBBBABABABABABABABAFEFEFFFFFFFFFFFFFF),
    .INIT_79(256'hFFFFFFFFFFFFFFFFFFBFBFBF96969696968686C6C6CEEFEFEFEDEDFDFDFDFDFD),
    .INIT_7A(256'hFDFDFDFDFDFDFD7F7F7F7F7F7F7F7F7FFFFFBFBABABABABABABAFAFAFEFFFFFF),
    .INIT_7B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFBFBFBF97969696968686C6C6CEEFEFEFEDEDFD),
    .INIT_7C(256'hEFEDEDFDFDFDFDFDFDFDFD7F7F7F7F7F7F7F7F7F7FBFBEBABABABABABABAFAFA),
    .INIT_7D(256'hBABAFAFAFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFBFB7969696968686C6C6C6CEEF),
    .INIT_7E(256'hC6C6CECFEFEDEDFDFDFDFDFDFDFDFDFF7F7F7F7F7F7F7F7F7FBFBEBEBABABABA),
    .INIT_7F(256'hBABABABABAFAFAFBFBFFFFFFFFFFFFFFFFFFFFFFFFFFBFBFB797969696868686),
    .MODE("SP16K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RSTBMUX("0"),
    .SRMODE("SYNC"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_5160x11_sub_000000_000 (
    .addra(addra[11:1]),
    .addrb(11'b00000000000),
    .bytea(addra[0]),
    .byteb(1'b0),
    .clka(clka),
    .csa(addra[12]),
    .dia({open_n51,open_n52,open_n53,open_n54,open_n55,open_n56,open_n57,open_n58,8'b00000000}),
    .rsta(rsta),
    .doa({open_n80,open_n81,open_n82,open_n83,open_n84,open_n85,open_n86,open_n87,inst_doa_i0_007,inst_doa_i0_006,inst_doa_i0_005,inst_doa_i0_004,inst_doa_i0_003,inst_doa_i0_002,inst_doa_i0_001,inst_doa_i0_000}));
  // address_offset=0;data_offset=8;depth=4096;width=3;num_section=1;width_per_section=3;section_size=11;working_depth=4096;working_width=8;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM32K #(
    .CLKBMUX("0"),
    .CSAMUX("INV"),
    .CSBMUX("0"),
    .DATA_WIDTH_A("8"),
    .DATA_WIDTH_B("8"),
    .INIT_00(256'h0707070707070707070707070707070707070707070707070707070707070707),
    .INIT_01(256'h0707070707070707070707070707070707070707070707070707070707070707),
    .INIT_02(256'h0707070707070707070707070707070707070707070707070707070707070707),
    .INIT_03(256'h0707070707070707070707070707070707070707070707070707070707070707),
    .INIT_04(256'h0707070707070707070707070707070707070707070707070707070707070707),
    .INIT_05(256'h0707070707070707070707070707070707070707070707070707070707070707),
    .INIT_06(256'h0707070707070707070707070707070707070707070707070707070707070707),
    .INIT_07(256'h0707070707070707070707070707070707070707070707070707070707070707),
    .INIT_08(256'h0707070707070707070707070707070404040404040707070707070707070707),
    .INIT_09(256'h0707070707070707070707070707070707070707070707070707070707070707),
    .INIT_0A(256'h0707070707070707070707070707040404040400000000000004040404040507),
    .INIT_0B(256'h0000000404070707070707070707070707070707070707070707070707070707),
    .INIT_0C(256'h0707070707070707070707070707070604000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000005070707070707070707070707070707070707070707),
    .INIT_0E(256'h0707070707070707070707070707070707060400000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000001070707070707070707070707070707),
    .INIT_10(256'h0707070707070707070707070707070707070707060000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000103070707070707070707),
    .INIT_12(256'h0707070707070707070707070707070707070707070707060000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000307070707),
    .INIT_14(256'h0707070707070707070707070707070707070707070707070706020000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000001),
    .INIT_16(256'h0000000005070707070707070707070707070707070707070707070707060000),
    .INIT_17(256'h0600000000000000000000000001030303030303030303020000000000000000),
    .INIT_18(256'h0000000000000000040507070707070707070707070707070707070707070707),
    .INIT_19(256'h0707070600000000000000000000000103030707070707070707070707020000),
    .INIT_1A(256'h0707060400000000000000000405070707070707070707070707070707070707),
    .INIT_1B(256'h0707070707070702000000000000000000000103070707070707070707070707),
    .INIT_1C(256'h0707070707070706040400000000000004040507070707070707070707070707),
    .INIT_1D(256'h0707070707070707070706000000000000000000000307070707070707070707),
    .INIT_1E(256'h0707070707070707070707070604040400000000040405050707070707070707),
    .INIT_1F(256'h0707070707070707070707070707020000000000000000000307070707070707),
    .INIT_20(256'h0707070707070707070707070707070707060404040000000404040507070707),
    .INIT_21(256'h0507070707070707070707070707070707060000000000000000000103070707),
    .INIT_22(256'h0707070707070707070707070707070707070707070606040404040004040405),
    .INIT_23(256'h0404040505070707070707070707070707070707070600000000000000000003),
    .INIT_24(256'h0000030707070707070707070707070707070707070707070707060404040404),
    .INIT_25(256'h0404040404040405050707070707070707070707070707070704000000000000),
    .INIT_26(256'h0000000000000307070707070707070707070707070707070707070707070606),
    .INIT_27(256'h0707060604040404040404040505070707070707070707070707070707040000),
    .INIT_28(256'h0400000000000000000203070707070707070707070707070707070707070707),
    .INIT_29(256'h0707070707070606040404040404040405050707070707070707070707070707),
    .INIT_2A(256'h0707070704000000000000000002070707070707070707070707070707070707),
    .INIT_2B(256'h0707070707070707070706060604040404040404050507070707070707070707),
    .INIT_2C(256'h0707070707070707040000000000000000020707070707070707070707070707),
    .INIT_2D(256'h0707070707070707070707070707060606040404040404040505070707070707),
    .INIT_2E(256'h0707070707070707070707070400000000000000020207070707070707070707),
    .INIT_2F(256'h0707070707070707070707070707070707070606060404040404040405050707),
    .INIT_30(256'h0505050707070707070707070707070504000000000000000202070707070707),
    .INIT_31(256'h0707070707070707070707070707070707070707070706060604040404040405),
    .INIT_32(256'h0404040505050507070707070707070707070705050400000000000002020707),
    .INIT_33(256'h0202030707070707070707070707070707070707070707070707060606040404),
    .INIT_34(256'h0604040404040405050505070707070707070707070707050504000000000000),
    .INIT_35(256'h0000000002020207070707070707070707070707070707070707070707060606),
    .INIT_36(256'h0706060606040404040405050505050707070707070707070707070505040000),
    .INIT_37(256'h0505000000000000020202070707070707070707070707070707070707070707),
    .INIT_38(256'h0707070706060606060404040404050505050507070707070707070707070705),
    .INIT_39(256'h0707070505050000000000000202020207070707070707070707070707070707),
    .INIT_3A(256'h0707070707070707060606060604040404050505050505070707070707070707),
    .INIT_3B(256'h0707070707070705050505000000000002020202070707070707070707070707),
    .INIT_3C(256'h0707070707070707070707060606060606040404040505050505050707070707),
    .INIT_3D(256'h0707070707070707070707050505050000000000020202020207070707070707),
    .INIT_3E(256'h0707070707070707070707070707060606060606060404040505050505050707),
    .INIT_3F(256'h0505070707070707070707070707070505050505000000000202020202060707),
    .INIT_40(256'h0202060607070707070707070707070706060606060606060404040505050505),
    .INIT_41(256'h0505050505050707070707070707070707070505050505050100000002020202),
    .INIT_42(256'h0202020202020206060607070707070707070606060606060606060604040505),
    .INIT_43(256'h0405050505050505050507070707070707070707070705050505050505000000),
    .INIT_44(256'h0505010000020202020202020606060606060606060606060606060606060606),
    .INIT_45(256'h0606060405050505050505050505070707070707070707070707050505050505),
    .INIT_46(256'h0505050505050501000202020202020202060606060606060606060606060606),
    .INIT_47(256'h0606060606060605050505050505050505070707070707070707070707070505),
    .INIT_48(256'h0707050505050505050505010100020202020202020206060606060606060606),
    .INIT_49(256'h0606060606060606060705050505050505050505050707070707070707070707),
    .INIT_4A(256'h0707070707070505050505050505050501010102020202020202020606060606),
    .INIT_4B(256'h0206060606060606060606060604050505050505050505050507070707070707),
    .INIT_4C(256'h0707070707070707070705050505050505050505050100020202020202020202),
    .INIT_4D(256'h0202020202020606060606060606060604040404050505050505050507070707),
    .INIT_4E(256'h0707070707070707070707070707050505050505050505050404000002020202),
    .INIT_4F(256'h0000020202020202020202060606060606060604040404040404050505050507),
    .INIT_50(256'h0505050707070707070707070707070707070505050505050505040404040404),
    .INIT_51(256'h0404040404000002020202020202020206060606060604040404040404040405),
    .INIT_52(256'h0404040405050707070707070707070707070707070705050505050505040404),
    .INIT_53(256'h0404040604040404040400000003030303030303030707040404040404040404),
    .INIT_54(256'h0404040404040404040707070707070707070707070707070707070505050505),
    .INIT_55(256'h0505050404040406060404040404040101010101010101010101050505040404),
    .INIT_56(256'h0505050404040404040404040406070707070707070707070707070707070705),
    .INIT_57(256'h0707070505050404040404060606040404050505010101010101010101010105),
    .INIT_58(256'h0101010505050505040404040404040606060607070707070707070707070707),
    .INIT_59(256'h0707070707070705050404040404040606060604050505050501010101010101),
    .INIT_5A(256'h0101010101010101050505050504040404040606060606070707070707070707),
    .INIT_5B(256'h0707070707070707070707050504040404040406060606070505050505050101),
    .INIT_5C(256'h0505050101010101010101010505050505050404040606060606060607070707),
    .INIT_5D(256'h0707070707070707070707070707070504040404040404060606070707050505),
    .INIT_5E(256'h0707050505050505010101010101010101050505050505060606060606060606),
    .INIT_5F(256'h0606060606070707070707070707070707070705040404040404040606070707),
    .INIT_60(256'h0607070707070707050505050101010101010101010505050507070606060606),
    .INIT_61(256'h0606060606060606060707070707070707070707070707040404040404040404),
    .INIT_62(256'h0404040407070707070707070707070705010101010101010107070707070707),
    .INIT_63(256'h0707070706060606060606060606070707070707070707070707070404040404),
    .INIT_64(256'h0404040404040404070707070707070707070707070303030303030303070707),
    .INIT_65(256'h0303070707070707070606060606060606060707070707070707070707070606),
    .INIT_66(256'h0707060604040404040404050707070707070707070707070703030303030303),
    .INIT_67(256'h0303030303030707070707070706060606060606060607070707070707070707),
    .INIT_68(256'h0707070707070606040404040404040507070707070707070707070707030303),
    .INIT_69(256'h0703030303030303030307070707070707060606060606060606070707070707),
    .INIT_6A(256'h0707070707070707070706060404040404040405050707070707070707070707),
    .INIT_6B(256'h0707070707030303030303030303070707070707070606060606060606060607),
    .INIT_6C(256'h0606060707070707070707070706060604040404040404050507070707070707),
    .INIT_6D(256'h0707070707070707070303030303030303030707070707070706060606060606),
    .INIT_6E(256'h0606060606060607070707070707070707060606060404040404040505070707),
    .INIT_6F(256'h0507070707070707070707070703030303030303030307070707070707060606),
    .INIT_70(256'h0706060606060606060606070707070707070707070606060604040404040405),
    .INIT_71(256'h0404040505050707070707070707070707030303030303030303070707070707),
    .INIT_72(256'h0707070707060606060606060606060707070707070707070706060606040404),
    .INIT_73(256'h0606040404040405050507070707070707070707070707070707070707070707),
    .INIT_74(256'h0707070707070707070606060606060606060607070707070707070707060606),
    .INIT_75(256'h0706060606060404040404050505050707070707070707070707070707070707),
    .INIT_76(256'h0707070707070707070707070706060606060606060607070707070707070707),
    .INIT_77(256'h0707070707070606060606040404040505050507070707070707070707070707),
    .INIT_78(256'h0707070707070707070707070707070706060606060606060606070707070707),
    .INIT_79(256'h0707070707070707070706060606060404040404050505050707070707070707),
    .INIT_7A(256'h0707070707070707070707070707070707070707060606060606060606060707),
    .INIT_7B(256'h0606070707070707070707070707060606060604040404040505050507070707),
    .INIT_7C(256'h0507070707070707070707070707070707070707070707070606060606060606),
    .INIT_7D(256'h0606060606070707070707070707070707070606060606060404040405050505),
    .INIT_7E(256'h0405050505050707070707070707070707070707070707070707070606060606),
    .INIT_7F(256'h0606060606060606060707070707070707070707070707060606060606040404),
    .MODE("SP16K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RSTBMUX("0"),
    .SRMODE("SYNC"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_5160x11_sub_000000_008 (
    .addra(addra[11:1]),
    .addrb(11'b00000000000),
    .bytea(addra[0]),
    .byteb(1'b0),
    .clka(clka),
    .csa(addra[12]),
    .dia({open_n108,open_n109,open_n110,open_n111,open_n112,open_n113,open_n114,open_n115,open_n116,open_n117,open_n118,open_n119,open_n120,3'b000}),
    .rsta(rsta),
    .doa({open_n142,open_n143,open_n144,open_n145,open_n146,open_n147,open_n148,open_n149,open_n150,open_n151,open_n152,open_n153,open_n154,inst_doa_i0_010,inst_doa_i0_009,inst_doa_i0_008}));
  // address_offset=4096;data_offset=0;depth=1064;width=11;num_section=1;width_per_section=11;section_size=11;working_depth=2048;working_width=16;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM32K #(
    .CLKBMUX("0"),
    .CSBMUX("0"),
    .DATA_WIDTH_A("16"),
    .DATA_WIDTH_B("16"),
    .INIT_00(256'h07FD07FD07FD07FF077F077F077F077F077F077F077F077F073F07BE06BE06BE),
    .INIT_01(256'h069604860486048604C604C605C605CE05EF05ED05ED07FD07FD07FD07FD07FD),
    .INIT_02(256'h07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07BF06BF06BF06B706960696),
    .INIT_03(256'h073E07BE06BE06BE06BA06BA06BA06BA06BA06FA06FA06F307FB07FF07FF07FF),
    .INIT_04(256'h07FD07FD07FD07FD07FD07FD07FD07FF077F077F077F077F077F077F077F073F),
    .INIT_05(256'h06BF06B7069706960696068604860486048604C604C605C605CF05ED05ED05FD),
    .INIT_06(256'h07FB07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF06BF),
    .INIT_07(256'h077F077F077F073F073E063E06BE06BE06BA06BA06BA06BA06FA06DA04F306F3),
    .INIT_08(256'h05CE05CD05ED05FD05FD07FD07FD07FD07FD07FD07FD07FF077F077F077F077F),
    .INIT_09(256'h07FF07FF07FF07BF06BF06BF06B7069606960686048604860486048604C604C6),
    .INIT_0A(256'h06D204D204F307F307FB07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF),
    .INIT_0B(256'h03FF037F037F037F037F077F073F073E063E063E06BE06BE06BA06BA06BA069A),
    .INIT_0C(256'h04860486048604C604C605C405CD05DD05FD05FD07FD07FD07FD07FD07FD03FF),
    .INIT_0D(256'h07FF07FF07FF07FF07FF07FF07FF07FF07BF06BF06B706970696068606860486),
    .INIT_0E(256'h06BA069A069A04D204D204D304F307F307FB07FF07FF07FF07FF07FF07FF07FF),
    .INIT_0F(256'h07FD07FD03FD03FF03FF037F037F037F037F033E063E063E063E063E06BE06BE),
    .INIT_10(256'h0697068606860686048604860486048604C604C405C405DC05DD05DD05FD05FD),
    .INIT_11(256'h07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07BF06BF06BF06B7),
    .INIT_12(256'h063A061A069A069A0492049204D204D204D304D305F307F307FB07FF07FF07FF),
    .INIT_13(256'h04D005D805D905D905F901F901F903FB03FB037B037B033A023A023A023A063A),
    .INIT_14(256'h07FB07BB06BB06BB06B30682068206820682048204820482048204C004C004D0),
    .INIT_15(256'h07FB07FB07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FB07FB),
    .INIT_16(256'h001A001A001A041A041A0412041204920492049204D204D204D305D305F307F3),
    .INIT_17(256'h04820480048004D004D004D004D004D804D800D800D800DA00DA001A001A001A),
    .INIT_18(256'h07FF07FF07FB07FB07FB07FB07BB06BB06B306A3068206820682068204820482),
    .INIT_19(256'h05D305D305F307F307FB07FB07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF),
    .INIT_1A(256'h009200120012001200120012001200120412041204120492049204D204D204D3),
    .INIT_1B(256'h0682068206820482048204800480049004900490049004900090009000900092),
    .INIT_1C(256'h07FF07FF07FF07FF07FF07FF07FB07FB07FB07FB07FB07BB06BB06A306A30682),
    .INIT_1D(256'h04D204D204D305D305D305D305F307F307FB07FB07FF07FF07FF07FF07FF07FF),
    .INIT_1E(256'h0090009000900092009200920012001200120012001200120412041204120492),
    .INIT_1F(256'h07BB06AB06A306A3068206820682068204820480048004900490049004900490),
    .INIT_20(256'h07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FB07FB07FB07FB07FB07FB),
    .INIT_21(256'h04120412041204D204D205D305D305D305D305D305F307F307FB07FB07FF07FF),
    .INIT_22(256'h0490049004900490009000900090009200920092001200120012001200120012),
    .INIT_23(256'h07FB07FB07FB07FB07FB07AB07AB06AB06A306A3068206820682068004800490),
    .INIT_24(256'h07FB07FB07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FB07FB),
    .INIT_25(256'h001200120012001204120412045204D305D305D305D305D305D305D305F307F3),
    .INIT_26(256'h0682068006800490049004900490049000900090009000920092009200120012),
    .INIT_27(256'h07FF07FF07FB07FB07FB07FB07FB07FB07FB07EB07AB07AB06AB06A306A30682),
    .INIT_28(256'h05D307F307FB07FB07FB07FB07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF),
    .INIT_29(256'h00920092001200120012001200120412045204530553055305D305D305D305D3),
    .INIT_2A(256'h07AB07AB06AB06A306A306A00680069006900690049004900490009000900092),
    .INIT_2B(256'h07FF07FF07FF07FF07FF07FF07FB07FB07FB07FB07FB07FB07FB07EB07EB07EB),
    .INIT_2C(256'h05D305D307F307F307FB07FB07FB07FB07FB07FB07FF07FF07FF07FF07FF07FF),
    .INIT_2D(256'h0490009000900092009200920012001200120012005205530553055305530553),
    .INIT_2E(256'h07FB07EB07EB07EB07EB07EB07AB07AB07AB06A106A106B00690069006900690),
    .INIT_2F(256'h07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FB07FB07FB07FB07FB07FB),
    .INIT_30(256'h057707770777077707F707FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF),
    .INIT_31(256'h07B507B507B506B506B406B40294029602960396019701170157015705570577),
    .INIT_32(256'h07FF07FF07FF07FF07FF07EF07EF07EF07EF07EF07EF07EF07AF07AD07AD07BD),
    .INIT_33(256'h07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF),
    .INIT_34(256'h07F707F707FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF),
    .INIT_35(256'h07FF07FF07FF07FF07FF07BF07BF07BF07BF07BF07BF07F703F703F703F703F7),
    .INIT_36(256'h07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF),
    .INIT_37(256'h07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF),
    .INIT_38(256'h07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF),
    .INIT_39(256'h07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF),
    .INIT_3A(256'h07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF),
    .INIT_3B(256'h07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF),
    .INIT_3C(256'h07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF),
    .INIT_3D(256'h07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF),
    .INIT_3E(256'h07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF),
    .INIT_3F(256'h07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF),
    .INIT_40(256'h07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF),
    .INIT_41(256'h07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF07FF),
    .INIT_42(256'h0000000000000000000000000000000007FF07FF07FF07FF07FF07FF07FF07FF),
    .INIT_43(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_44(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_45(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_46(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_47(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_48(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_49(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_50(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_51(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_52(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_53(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_54(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_55(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_56(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_57(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_58(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_59(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_60(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_61(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_62(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_63(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_64(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_65(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_66(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_67(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_68(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_69(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_70(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_71(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_72(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_73(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_74(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_75(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_76(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_77(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_78(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_79(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP16K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RSTBMUX("0"),
    .SRMODE("SYNC"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_5160x11_sub_004096_000 (
    .addra(addra[10:0]),
    .addrb(11'b00000000000),
    .bytewea(1'b0),
    .byteweb(1'b0),
    .clka(clka),
    .csa(\and_Naddra[11]_addra_o ),
    .dia({open_n175,open_n176,open_n177,open_n178,open_n179,11'b00000000000}),
    .rsta(rsta),
    .doa({open_n201,open_n202,open_n203,open_n204,open_n205,inst_doa_i2_010,inst_doa_i2_009,inst_doa_i2_008,inst_doa_i2_007,inst_doa_i2_006,inst_doa_i2_005,inst_doa_i2_004,inst_doa_i2_003,inst_doa_i2_002,inst_doa_i2_001,inst_doa_i2_000}));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_0  (
    .i0(inst_doa_i0_000),
    .i1(inst_doa_i0_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_0 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_1  (
    .i0(inst_doa_i2_000),
    .i1(inst_doa_i2_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_1 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b0/B0_0 ),
    .i1(\inst_doa_mux_b0/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[0]));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_0  (
    .i0(inst_doa_i0_001),
    .i1(inst_doa_i0_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_0 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_1  (
    .i0(inst_doa_i2_001),
    .i1(inst_doa_i2_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_1 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b1/B0_0 ),
    .i1(\inst_doa_mux_b1/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[1]));
  AL_MUX \inst_doa_mux_b10/al_mux_b0_0_0  (
    .i0(inst_doa_i0_010),
    .i1(inst_doa_i0_010),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b10/B0_0 ));
  AL_MUX \inst_doa_mux_b10/al_mux_b0_0_1  (
    .i0(inst_doa_i2_010),
    .i1(inst_doa_i2_010),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b10/B0_1 ));
  AL_MUX \inst_doa_mux_b10/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b10/B0_0 ),
    .i1(\inst_doa_mux_b10/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[10]));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_0  (
    .i0(inst_doa_i0_002),
    .i1(inst_doa_i0_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_0 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_1  (
    .i0(inst_doa_i2_002),
    .i1(inst_doa_i2_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_1 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b2/B0_0 ),
    .i1(\inst_doa_mux_b2/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[2]));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_0  (
    .i0(inst_doa_i0_003),
    .i1(inst_doa_i0_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_0 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_1  (
    .i0(inst_doa_i2_003),
    .i1(inst_doa_i2_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_1 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b3/B0_0 ),
    .i1(\inst_doa_mux_b3/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[3]));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_0  (
    .i0(inst_doa_i0_004),
    .i1(inst_doa_i0_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_0 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_1  (
    .i0(inst_doa_i2_004),
    .i1(inst_doa_i2_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_1 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b4/B0_0 ),
    .i1(\inst_doa_mux_b4/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[4]));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_0  (
    .i0(inst_doa_i0_005),
    .i1(inst_doa_i0_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_0 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_1  (
    .i0(inst_doa_i2_005),
    .i1(inst_doa_i2_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_1 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b5/B0_0 ),
    .i1(\inst_doa_mux_b5/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[5]));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_0  (
    .i0(inst_doa_i0_006),
    .i1(inst_doa_i0_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_0 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_1  (
    .i0(inst_doa_i2_006),
    .i1(inst_doa_i2_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_1 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b6/B0_0 ),
    .i1(\inst_doa_mux_b6/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[6]));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_0  (
    .i0(inst_doa_i0_007),
    .i1(inst_doa_i0_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_0 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_1  (
    .i0(inst_doa_i2_007),
    .i1(inst_doa_i2_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_1 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b7/B0_0 ),
    .i1(\inst_doa_mux_b7/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[7]));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_0  (
    .i0(inst_doa_i0_008),
    .i1(inst_doa_i0_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_0 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_1  (
    .i0(inst_doa_i2_008),
    .i1(inst_doa_i2_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_1 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b8/B0_0 ),
    .i1(\inst_doa_mux_b8/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[8]));
  AL_MUX \inst_doa_mux_b9/al_mux_b0_0_0  (
    .i0(inst_doa_i0_009),
    .i1(inst_doa_i0_009),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b9/B0_0 ));
  AL_MUX \inst_doa_mux_b9/al_mux_b0_0_1  (
    .i0(inst_doa_i2_009),
    .i1(inst_doa_i2_009),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b9/B0_1 ));
  AL_MUX \inst_doa_mux_b9/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b9/B0_0 ),
    .i1(\inst_doa_mux_b9/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[9]));

endmodule 

