// Verilog netlist created by TD v4.6.18154
// Fri Nov 13 11:12:27 2020

`timescale 1ns / 1ps
module its  // al_ip/word/its.v(14)
  (
  addra,
  clka,
  rsta,
  doa
  );

  input [13:0] addra;  // al_ip/word/its.v(18)
  input clka;  // al_ip/word/its.v(19)
  input rsta;  // al_ip/word/its.v(20)
  output [0:0] doa;  // al_ip/word/its.v(16)

  wire [0:0] addra_piped;
  wire inst_doa_i0_000;
  wire inst_doa_i1_000;

  reg_sr_as_w1 addra_pipe (
    .clk(clka),
    .d(addra[13]),
    .en(1'b1),
    .reset(rsta),
    .set(1'b0),
    .q(addra_piped));
  EG_PHY_CONFIG #(
    .DONE_PERSISTN("ENABLE"),
    .INIT_PERSISTN("ENABLE"),
    .JTAG_PERSISTN("DISABLE"),
    .PROGRAMN_PERSISTN("DISABLE"))
    config_inst ();
  // address_offset=0;data_offset=0;depth=8192;width=1;num_section=1;width_per_section=1;section_size=1;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_02(256'hFFFFFFF803FFFFFFFFFFFFF801FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_03(256'hFFFFF803FFFFFFFFFFFFF801FFFFFFFFFFFFFF803FFFFFFFFFFFFF801FFFFFFF),
    .INIT_04(256'hFFF803FFFFFFFFFFFFF801FFFFFFFFFFFFFF803FFFFFFFFFFFFF801FFFFFFFFF),
    .INIT_05(256'hF803FFFFFDFFFFFFF801FFFFFFFFFFFFFF803FFFFFFFFFFFFF801FFFFFFFFFFF),
    .INIT_06(256'h03FFFFFC07FFFFF801FFFFFFFFFFFFFF803FFFFFC3FFFFFF801FFFFFFFFFFFFF),
    .INIT_07(256'hFFFFFC00FFFFF801FFFFFFFFFFFFFF803FFFFFC00FFFFF801FFFFFFFFFFFFFF8),
    .INIT_08(256'hFFFC00FFFFF801FFFFFFFFFFFFFFC07FFFFFC00FFFFF801FFFFFFFFFFFFFF803),
    .INIT_09(256'hFC00FFFFF801FFFFFFFFFFFFFFC07FFFFFC00FFFFF801FFFFFFFFFFFFFFC07FF),
    .INIT_0A(256'h00FFFFF801FFFFFFFFFFFFFFC07FFFFFC00FFFFF801FFFFFFFFFFFFFFC07FFFF),
    .INIT_0B(256'hFFFFF801FFFFFFFFFFFFFFC07FFFFFC00FFFFF801FFFFFFFFFFFFFFC07FFFFFC),
    .INIT_0C(256'hFFF801FFFFFFFFFFFFFFC07FFFFFC00FFFFF801FFFFFFFFFFFFFFC07FFFFFC00),
    .INIT_0D(256'hF801FFFFE03FFFFFFFC07FFFFFC00FFFFF801FFFFFFFFFFFFFFC07FFFFFC00FF),
    .INIT_0E(256'h01FFE000007FFFFFC07FFC00000007FF801FFFC0001FFFFFFC07FFC00000007F),
    .INIT_0F(256'hFFC0000007FFFFFFFFFC00000007FF801FFC000001FFFFFFFFFFC00000007FF8),
    .INIT_10(256'hC0000001FFFFFFFFFC00000007FF801FFC0000003FFFFFFFFFC00000007FF801),
    .INIT_11(256'hFFF8007FFFFFFFFC00000007FF801FFC0078000FFFFFFFFFC00000007FF801FF),
    .INIT_12(256'hFE003FFFFFFFFFFFC00FFFFF801FFC3FFFC007FFFFFFFFFFFC00FFFFF801FFC0),
    .INIT_13(256'h803FFFFFFFFFFFC00FFFFF801FFFFFFFF003FFFFFFFFFFFC00FFFFF801FFCFFF),
    .INIT_14(256'h1FFFFFFFFFFFC00FFFFF801FFFFFFFF801FFFFFFFFFFFC00FFFFF801FFFFFFFF),
    .INIT_15(256'hFFFFFFFFFFC00FFFFF801FFFFFFFF801FFFFFFFFFFFC00FFFFF801FFFFFFFF80),
    .INIT_16(256'hFFFFFFFFC00FFFFF801FFFFFFFF801FFFFFFFFFFFC00FFFFF801FFFFFFFF801F),
    .INIT_17(256'hFFFFFFC00FFFFF801FFFFFFFF003FFFFFFFFFFFC00FFFFF801FFFFFFFF003FFF),
    .INIT_18(256'hFFFFC00FFFFF801FFFFFFF8003FFFFFFFFFFFC00FFFFF801FFFFFFFC003FFFFF),
    .INIT_19(256'hFFC00FFFFF801FFFFFF80007FFFFFFFFFFFC00FFFFF801FFFFFFE0007FFFFFFF),
    .INIT_1A(256'hC00FFFFF801FFFFF00001FFFFFFFFFFFFC00FFFFF801FFFFFC0000FFFFFFFFFF),
    .INIT_1B(256'h0FFFFF801FFFF00000FFFFFFFFFFFFFC00FFFFF801FFFFC00003FFFFFFFFFFFF),
    .INIT_1C(256'hFFFF801FFF00000FFFFFFFFFFFFFFC00FFFFF801FFFC00003FFFFFFFFFFFFFC0),
    .INIT_1D(256'hFF801FFC0000FFFFFFFFFFFFFFFC00FFFFF801FFE00003FFFFFFFFFFFFFFC00F),
    .INIT_1E(256'h801FF8001FFFFFFFFFFFFFFFFC00FFFFF801FF80007FFFFFFFFFFFFFFFC00FFF),
    .INIT_1F(256'h1FF000FFFFFFFFFFFFFFFFFC00FFFFF801FF0007FFFFFFFFFFFFFFFFC00FFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_11352x1_sub_000000_000 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n63,open_n64,addra[13]}),
    .dia({open_n68,open_n69,open_n70,open_n71,open_n72,open_n73,open_n74,1'b0,open_n75}),
    .rsta(rsta),
    .doa({open_n90,open_n91,open_n92,open_n93,open_n94,open_n95,open_n96,open_n97,inst_doa_i0_000}));
  // address_offset=8192;data_offset=0;depth=3160;width=1;num_section=1;width_per_section=1;section_size=1;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hF003FFFFFFFFFFFFFFFFFC00FFFFF801FF001FFFFFFFFFFFFFFFFFC00FFFFF80),
    .INIT_01(256'h07FFFFFFFFFFFFFFFFFC00FFFFF801FE007FFFFFFFFFFFFFFFFFC00FFFFF801F),
    .INIT_02(256'hFFFFFFFFFFFFFFFFFC00FFFFF801FE007FFFFFFFFFFFFFFFFFC00FFFFF801FE0),
    .INIT_03(256'hFFFFFFFFFFFFFFFC01FFFFF801FE007FFFFFFFFFFFFFFFFFC00FFFFF801FE007),
    .INIT_04(256'hF1FFFFFFFFFFF801FFFFF801FF003FFFFF9FFFFFFFFFFF801FFFFF801FF007FF),
    .INIT_05(256'hFFFFFFFFCFE001FFFFF801FF801FFFFC1FFFFFFFFFFF001FFFFF801FF003FFFF),
    .INIT_06(256'hFFFFFFC00003FFFFF801FFC0007C001FFFFFFFFC00003FFFFF801FF8007FFE01),
    .INIT_07(256'hFFFFC00007FFFFF801FFF00000001FFFFFFFFC00007FFFFF801FFE00000001FF),
    .INIT_08(256'hFFC0001FFFFFF801FFFE0000001FFFFFFFFC0000FFFFFF801FFF80000001FFFF),
    .INIT_09(256'hFE07FFFFFFFFFFFFFFE00003FFFFFFFFFF0007FFFFFF801FFFF8000007FFFFFF),
    .INIT_0A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80FFFFFFFFFFF),
    .INIT_0B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0C(256'h000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_11352x1_sub_008192_000 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n123,open_n124,addra[13]}),
    .dia({open_n128,open_n129,open_n130,open_n131,open_n132,open_n133,open_n134,1'b0,open_n135}),
    .rsta(rsta),
    .doa({open_n150,open_n151,open_n152,open_n153,open_n154,open_n155,open_n156,open_n157,inst_doa_i1_000}));
  AL_MUX \inst_doa_mux/al_mux_b0_0_0  (
    .i0(inst_doa_i0_000),
    .i1(inst_doa_i1_000),
    .sel(addra_piped),
    .o(doa));

endmodule 

